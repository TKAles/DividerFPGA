-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Aug 2 2023 08:20:12

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    sr_sel_row : in std_logic;
    sr_sel_div : in std_logic;
    sr_clk : in std_logic;
    row_completed : out std_logic;
    en_internals : in std_logic;
    divide_enable : in std_logic;
    sr_reset : in std_logic;
    laser_pulse : in std_logic;
    sr_data : in std_logic;
    en_rowpack : in std_logic;
    divided_pulse : out std_logic;
    constant_v : in std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__5170\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4248\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4219\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4186\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4120\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4054\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4030\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4008\ : std_logic;
signal \N__4005\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3993\ : std_logic;
signal \N__3990\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3984\ : std_logic;
signal \N__3981\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3975\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3963\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3919\ : std_logic;
signal \N__3916\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3910\ : std_logic;
signal \N__3907\ : std_logic;
signal \N__3904\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3894\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3886\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3879\ : std_logic;
signal \N__3878\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3867\ : std_logic;
signal \N__3862\ : std_logic;
signal \N__3859\ : std_logic;
signal \N__3856\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3846\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3821\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3817\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3799\ : std_logic;
signal \N__3796\ : std_logic;
signal \N__3793\ : std_logic;
signal \N__3790\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3771\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3756\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3744\ : std_logic;
signal \N__3741\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3726\ : std_logic;
signal \N__3723\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3711\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3696\ : std_logic;
signal \N__3693\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3681\ : std_logic;
signal \N__3678\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3663\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3651\ : std_logic;
signal \N__3648\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3633\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3620\ : std_logic;
signal \N__3617\ : std_logic;
signal \N__3614\ : std_logic;
signal \N__3609\ : std_logic;
signal \N__3606\ : std_logic;
signal \N__3603\ : std_logic;
signal \N__3600\ : std_logic;
signal \N__3597\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3593\ : std_logic;
signal \N__3590\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3582\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3573\ : std_logic;
signal \N__3572\ : std_logic;
signal \N__3569\ : std_logic;
signal \N__3566\ : std_logic;
signal \N__3561\ : std_logic;
signal \N__3558\ : std_logic;
signal \N__3555\ : std_logic;
signal \N__3552\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3548\ : std_logic;
signal \N__3545\ : std_logic;
signal \N__3540\ : std_logic;
signal \N__3537\ : std_logic;
signal \N__3536\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3530\ : std_logic;
signal \N__3525\ : std_logic;
signal \N__3522\ : std_logic;
signal \N__3519\ : std_logic;
signal \N__3516\ : std_logic;
signal \N__3513\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3501\ : std_logic;
signal \N__3498\ : std_logic;
signal \N__3497\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3491\ : std_logic;
signal \N__3486\ : std_logic;
signal \N__3483\ : std_logic;
signal \N__3482\ : std_logic;
signal \N__3479\ : std_logic;
signal \N__3476\ : std_logic;
signal \N__3471\ : std_logic;
signal \N__3468\ : std_logic;
signal \N__3465\ : std_logic;
signal \N__3462\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3456\ : std_logic;
signal \N__3453\ : std_logic;
signal \N__3450\ : std_logic;
signal \N__3447\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3441\ : std_logic;
signal \N__3438\ : std_logic;
signal \N__3437\ : std_logic;
signal \N__3434\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3428\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3417\ : std_logic;
signal \N__3416\ : std_logic;
signal \N__3413\ : std_logic;
signal \N__3410\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3402\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3396\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3390\ : std_logic;
signal \N__3389\ : std_logic;
signal \N__3388\ : std_logic;
signal \N__3385\ : std_logic;
signal \N__3380\ : std_logic;
signal \N__3375\ : std_logic;
signal \N__3374\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3368\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3361\ : std_logic;
signal \N__3358\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3350\ : std_logic;
signal \N__3347\ : std_logic;
signal \N__3344\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3334\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3324\ : std_logic;
signal \N__3321\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3319\ : std_logic;
signal \N__3318\ : std_logic;
signal \N__3317\ : std_logic;
signal \N__3316\ : std_logic;
signal \N__3315\ : std_logic;
signal \N__3312\ : std_logic;
signal \N__3303\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3298\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3295\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3290\ : std_logic;
signal \N__3289\ : std_logic;
signal \N__3286\ : std_logic;
signal \N__3283\ : std_logic;
signal \N__3270\ : std_logic;
signal \N__3261\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3248\ : std_logic;
signal \N__3245\ : std_logic;
signal \N__3244\ : std_logic;
signal \N__3243\ : std_logic;
signal \N__3242\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3238\ : std_logic;
signal \N__3237\ : std_logic;
signal \N__3236\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3228\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3222\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3220\ : std_logic;
signal \N__3217\ : std_logic;
signal \N__3216\ : std_logic;
signal \N__3213\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3211\ : std_logic;
signal \N__3210\ : std_logic;
signal \N__3207\ : std_logic;
signal \N__3204\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3186\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3176\ : std_logic;
signal \N__3165\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3160\ : std_logic;
signal \N__3157\ : std_logic;
signal \N__3154\ : std_logic;
signal \N__3151\ : std_logic;
signal \N__3148\ : std_logic;
signal \N__3141\ : std_logic;
signal \N__3140\ : std_logic;
signal \N__3137\ : std_logic;
signal \N__3134\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3121\ : std_logic;
signal \N__3114\ : std_logic;
signal \N__3111\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3109\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3103\ : std_logic;
signal \N__3100\ : std_logic;
signal \N__3093\ : std_logic;
signal \N__3090\ : std_logic;
signal \N__3087\ : std_logic;
signal \N__3084\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3078\ : std_logic;
signal \N__3075\ : std_logic;
signal \N__3072\ : std_logic;
signal \N__3069\ : std_logic;
signal \N__3066\ : std_logic;
signal \N__3063\ : std_logic;
signal \N__3060\ : std_logic;
signal \N__3057\ : std_logic;
signal \N__3054\ : std_logic;
signal \N__3051\ : std_logic;
signal \N__3048\ : std_logic;
signal \N__3047\ : std_logic;
signal \N__3044\ : std_logic;
signal \N__3043\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3037\ : std_logic;
signal \N__3034\ : std_logic;
signal \N__3027\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3022\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3012\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3010\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3002\ : std_logic;
signal \N__2997\ : std_logic;
signal \N__2996\ : std_logic;
signal \N__2993\ : std_logic;
signal \N__2992\ : std_logic;
signal \N__2989\ : std_logic;
signal \N__2986\ : std_logic;
signal \N__2983\ : std_logic;
signal \N__2976\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2974\ : std_logic;
signal \N__2971\ : std_logic;
signal \N__2968\ : std_logic;
signal \N__2965\ : std_logic;
signal \N__2958\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2956\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2948\ : std_logic;
signal \N__2943\ : std_logic;
signal \N__2942\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2938\ : std_logic;
signal \N__2933\ : std_logic;
signal \N__2928\ : std_logic;
signal \N__2927\ : std_logic;
signal \N__2924\ : std_logic;
signal \N__2923\ : std_logic;
signal \N__2920\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2914\ : std_logic;
signal \N__2907\ : std_logic;
signal \N__2904\ : std_logic;
signal \N__2901\ : std_logic;
signal \N__2898\ : std_logic;
signal \N__2895\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2889\ : std_logic;
signal \N__2886\ : std_logic;
signal \N__2883\ : std_logic;
signal \N__2880\ : std_logic;
signal \N__2877\ : std_logic;
signal \N__2876\ : std_logic;
signal \N__2871\ : std_logic;
signal \N__2868\ : std_logic;
signal \N__2865\ : std_logic;
signal \N__2862\ : std_logic;
signal \N__2859\ : std_logic;
signal \N__2856\ : std_logic;
signal \N__2855\ : std_logic;
signal \N__2850\ : std_logic;
signal \N__2847\ : std_logic;
signal \N__2844\ : std_logic;
signal \N__2841\ : std_logic;
signal \N__2838\ : std_logic;
signal \N__2837\ : std_logic;
signal \N__2836\ : std_logic;
signal \N__2835\ : std_logic;
signal \N__2830\ : std_logic;
signal \N__2825\ : std_logic;
signal \N__2820\ : std_logic;
signal \N__2817\ : std_logic;
signal \N__2814\ : std_logic;
signal \N__2811\ : std_logic;
signal \N__2808\ : std_logic;
signal \N__2807\ : std_logic;
signal \N__2806\ : std_logic;
signal \N__2803\ : std_logic;
signal \N__2798\ : std_logic;
signal \N__2793\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2781\ : std_logic;
signal \N__2780\ : std_logic;
signal \N__2779\ : std_logic;
signal \N__2776\ : std_logic;
signal \N__2771\ : std_logic;
signal \N__2766\ : std_logic;
signal \N__2763\ : std_logic;
signal \N__2760\ : std_logic;
signal \N__2757\ : std_logic;
signal \N__2754\ : std_logic;
signal \N__2751\ : std_logic;
signal \N__2748\ : std_logic;
signal \N__2745\ : std_logic;
signal \N__2742\ : std_logic;
signal \N__2739\ : std_logic;
signal \N__2736\ : std_logic;
signal \N__2733\ : std_logic;
signal \N__2730\ : std_logic;
signal \N__2727\ : std_logic;
signal \N__2724\ : std_logic;
signal \N__2721\ : std_logic;
signal \N__2718\ : std_logic;
signal \N__2715\ : std_logic;
signal \N__2712\ : std_logic;
signal \N__2709\ : std_logic;
signal \N__2706\ : std_logic;
signal \N__2703\ : std_logic;
signal \N__2700\ : std_logic;
signal \N__2697\ : std_logic;
signal \N__2694\ : std_logic;
signal \N__2691\ : std_logic;
signal \N__2688\ : std_logic;
signal \N__2685\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2679\ : std_logic;
signal \N__2676\ : std_logic;
signal \N__2673\ : std_logic;
signal \N__2670\ : std_logic;
signal \N__2667\ : std_logic;
signal \N__2664\ : std_logic;
signal \N__2661\ : std_logic;
signal \N__2658\ : std_logic;
signal \N__2655\ : std_logic;
signal \N__2652\ : std_logic;
signal \N__2649\ : std_logic;
signal \N__2648\ : std_logic;
signal \N__2647\ : std_logic;
signal \N__2646\ : std_logic;
signal \N__2641\ : std_logic;
signal \N__2636\ : std_logic;
signal \N__2631\ : std_logic;
signal \N__2630\ : std_logic;
signal \N__2629\ : std_logic;
signal \N__2628\ : std_logic;
signal \N__2619\ : std_logic;
signal \N__2616\ : std_logic;
signal \N__2613\ : std_logic;
signal \N__2610\ : std_logic;
signal \N__2607\ : std_logic;
signal \N__2604\ : std_logic;
signal \N__2601\ : std_logic;
signal \N__2598\ : std_logic;
signal \N__2595\ : std_logic;
signal \N__2592\ : std_logic;
signal \N__2589\ : std_logic;
signal \N__2586\ : std_logic;
signal \N__2583\ : std_logic;
signal \N__2580\ : std_logic;
signal \N__2577\ : std_logic;
signal \N__2574\ : std_logic;
signal \N__2571\ : std_logic;
signal \N__2568\ : std_logic;
signal \N__2565\ : std_logic;
signal \N__2562\ : std_logic;
signal \N__2559\ : std_logic;
signal \N__2556\ : std_logic;
signal \N__2553\ : std_logic;
signal \N__2550\ : std_logic;
signal \N__2547\ : std_logic;
signal \N__2544\ : std_logic;
signal \N__2541\ : std_logic;
signal \N__2540\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2534\ : std_logic;
signal \N__2531\ : std_logic;
signal \N__2526\ : std_logic;
signal \N__2523\ : std_logic;
signal \N__2522\ : std_logic;
signal \N__2519\ : std_logic;
signal \N__2516\ : std_logic;
signal \N__2513\ : std_logic;
signal \N__2508\ : std_logic;
signal \N__2505\ : std_logic;
signal \N__2502\ : std_logic;
signal \N__2499\ : std_logic;
signal \N__2496\ : std_logic;
signal \N__2493\ : std_logic;
signal \N__2490\ : std_logic;
signal \N__2487\ : std_logic;
signal \N__2484\ : std_logic;
signal \N__2481\ : std_logic;
signal \N__2478\ : std_logic;
signal \N__2475\ : std_logic;
signal \N__2472\ : std_logic;
signal \N__2469\ : std_logic;
signal \N__2466\ : std_logic;
signal \N__2463\ : std_logic;
signal \N__2460\ : std_logic;
signal \N__2457\ : std_logic;
signal \N__2454\ : std_logic;
signal \N__2451\ : std_logic;
signal \N__2448\ : std_logic;
signal \N__2445\ : std_logic;
signal \N__2442\ : std_logic;
signal \N__2439\ : std_logic;
signal \N__2436\ : std_logic;
signal \N__2433\ : std_logic;
signal \N__2430\ : std_logic;
signal \N__2427\ : std_logic;
signal \N__2424\ : std_logic;
signal \N__2421\ : std_logic;
signal \N__2420\ : std_logic;
signal \N__2417\ : std_logic;
signal \N__2414\ : std_logic;
signal \N__2409\ : std_logic;
signal \N__2406\ : std_logic;
signal \N__2405\ : std_logic;
signal \N__2402\ : std_logic;
signal \N__2399\ : std_logic;
signal \N__2394\ : std_logic;
signal \N__2391\ : std_logic;
signal \N__2390\ : std_logic;
signal \N__2387\ : std_logic;
signal \N__2384\ : std_logic;
signal \N__2379\ : std_logic;
signal \N__2376\ : std_logic;
signal \N__2375\ : std_logic;
signal \N__2372\ : std_logic;
signal \N__2369\ : std_logic;
signal \N__2364\ : std_logic;
signal \N__2361\ : std_logic;
signal \N__2360\ : std_logic;
signal \N__2357\ : std_logic;
signal \N__2354\ : std_logic;
signal \N__2349\ : std_logic;
signal \N__2346\ : std_logic;
signal \N__2345\ : std_logic;
signal \N__2342\ : std_logic;
signal \N__2339\ : std_logic;
signal \N__2334\ : std_logic;
signal \N__2331\ : std_logic;
signal \N__2330\ : std_logic;
signal \N__2327\ : std_logic;
signal \N__2324\ : std_logic;
signal \N__2319\ : std_logic;
signal \N__2316\ : std_logic;
signal \N__2315\ : std_logic;
signal \N__2312\ : std_logic;
signal \N__2309\ : std_logic;
signal \N__2304\ : std_logic;
signal \N__2301\ : std_logic;
signal \N__2300\ : std_logic;
signal \N__2297\ : std_logic;
signal \N__2294\ : std_logic;
signal \N__2289\ : std_logic;
signal \N__2286\ : std_logic;
signal \N__2283\ : std_logic;
signal \N__2282\ : std_logic;
signal \N__2277\ : std_logic;
signal \N__2274\ : std_logic;
signal \N__2271\ : std_logic;
signal \N__2268\ : std_logic;
signal \N__2265\ : std_logic;
signal \N__2262\ : std_logic;
signal \N__2261\ : std_logic;
signal \N__2258\ : std_logic;
signal \N__2255\ : std_logic;
signal \N__2250\ : std_logic;
signal \N__2247\ : std_logic;
signal \N__2244\ : std_logic;
signal \N__2243\ : std_logic;
signal \N__2240\ : std_logic;
signal \N__2237\ : std_logic;
signal \N__2232\ : std_logic;
signal \N__2229\ : std_logic;
signal \N__2226\ : std_logic;
signal \N__2223\ : std_logic;
signal \N__2220\ : std_logic;
signal \N__2217\ : std_logic;
signal \N__2214\ : std_logic;
signal \N__2213\ : std_logic;
signal \N__2210\ : std_logic;
signal \N__2207\ : std_logic;
signal \N__2202\ : std_logic;
signal \N__2199\ : std_logic;
signal \N__2198\ : std_logic;
signal \N__2195\ : std_logic;
signal \N__2192\ : std_logic;
signal \N__2187\ : std_logic;
signal \N__2184\ : std_logic;
signal \N__2183\ : std_logic;
signal \N__2180\ : std_logic;
signal \N__2177\ : std_logic;
signal \N__2172\ : std_logic;
signal \N__2169\ : std_logic;
signal \N__2168\ : std_logic;
signal \N__2165\ : std_logic;
signal \N__2162\ : std_logic;
signal \N__2157\ : std_logic;
signal \N__2154\ : std_logic;
signal \N__2153\ : std_logic;
signal \N__2150\ : std_logic;
signal \N__2147\ : std_logic;
signal \N__2142\ : std_logic;
signal \N__2139\ : std_logic;
signal \N__2136\ : std_logic;
signal \N__2133\ : std_logic;
signal \N__2130\ : std_logic;
signal \N__2127\ : std_logic;
signal \N__2124\ : std_logic;
signal \N__2121\ : std_logic;
signal \N__2118\ : std_logic;
signal \N__2115\ : std_logic;
signal \N__2112\ : std_logic;
signal \N__2109\ : std_logic;
signal \N__2106\ : std_logic;
signal \N__2103\ : std_logic;
signal \N__2100\ : std_logic;
signal \N__2097\ : std_logic;
signal \N__2094\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \bfn_1_7_0_\ : std_logic;
signal \pulse_counter.n728\ : std_logic;
signal \pulse_counter.n729\ : std_logic;
signal \pulse_counter.n730\ : std_logic;
signal \pulse_counter.n731\ : std_logic;
signal \pulse_counter.n732\ : std_logic;
signal \pulse_counter.n733\ : std_logic;
signal \pulse_counter.n734\ : std_logic;
signal \pulse_counter.n735\ : std_logic;
signal \bfn_1_8_0_\ : std_logic;
signal \pulse_counter.n736\ : std_logic;
signal \pulse_counter.n737\ : std_logic;
signal \pulse_counter.n738\ : std_logic;
signal \pulse_counter.n739\ : std_logic;
signal \pulse_counter.n740\ : std_logic;
signal \pulse_counter.n741\ : std_logic;
signal \pulse_counter.n742\ : std_logic;
signal divide_enable_c : std_logic;
signal n176 : std_logic;
signal output_state : std_logic;
signal constant_v_c : std_logic;
signal \pulse_counter.internal_count_0\ : std_logic;
signal \bfn_2_7_0_\ : std_logic;
signal \pulse_counter.internal_count_1\ : std_logic;
signal \pulse_counter.n712\ : std_logic;
signal \pulse_counter.internal_count_2\ : std_logic;
signal \pulse_counter.n713\ : std_logic;
signal \pulse_counter.internal_count_3\ : std_logic;
signal \pulse_counter.n714\ : std_logic;
signal \pulse_counter.internal_count_4\ : std_logic;
signal \pulse_counter.n715\ : std_logic;
signal \pulse_counter.internal_count_5\ : std_logic;
signal \pulse_counter.n716\ : std_logic;
signal \pulse_counter.internal_count_6\ : std_logic;
signal \pulse_counter.n717\ : std_logic;
signal \pulse_counter.internal_count_7\ : std_logic;
signal \pulse_counter.n718\ : std_logic;
signal \pulse_counter.n719\ : std_logic;
signal \pulse_counter.internal_count_8\ : std_logic;
signal \bfn_2_8_0_\ : std_logic;
signal \pulse_counter.internal_count_9\ : std_logic;
signal \pulse_counter.n720\ : std_logic;
signal \pulse_counter.internal_count_10\ : std_logic;
signal \pulse_counter.n721\ : std_logic;
signal \pulse_counter.internal_count_11\ : std_logic;
signal \pulse_counter.n722\ : std_logic;
signal \pulse_counter.internal_count_12\ : std_logic;
signal \pulse_counter.n723\ : std_logic;
signal \pulse_counter.internal_count_13\ : std_logic;
signal \pulse_counter.n724\ : std_logic;
signal \pulse_counter.internal_count_14\ : std_logic;
signal \pulse_counter.n725\ : std_logic;
signal \pulse_counter.internal_count_15\ : std_logic;
signal \pulse_counter.n726\ : std_logic;
signal \pulse_counter.n727\ : std_logic;
signal \pulse_counter.n13\ : std_logic;
signal \bfn_2_9_0_\ : std_logic;
signal n4_adj_116 : std_logic;
signal n5_adj_120 : std_logic;
signal n1_adj_117 : std_logic;
signal n9 : std_logic;
signal \n795_cascade_\ : std_logic;
signal n6_adj_119 : std_logic;
signal n12 : std_logic;
signal n16 : std_logic;
signal \n817_cascade_\ : std_logic;
signal n787 : std_logic;
signal \n825_cascade_\ : std_logic;
signal sr_divider_data_11 : std_logic;
signal sr_divider_data_13 : std_logic;
signal count_done : std_logic;
signal laser_pulse_c : std_logic;
signal sr_divider_data_2 : std_logic;
signal sr_divider_data_14 : std_logic;
signal sr_divider_data_15 : std_logic;
signal sr_divider_data_0 : std_logic;
signal sr_divider_data_3 : std_logic;
signal sr_divider_data_12 : std_logic;
signal sr_divider_data_1 : std_logic;
signal sr_divider_data_10 : std_logic;
signal sr_divider_data_6 : std_logic;
signal sr_divider_data_9 : std_logic;
signal sr_divider_data_4 : std_logic;
signal sr_divider_data_5 : std_logic;
signal sr_divider_data_8 : std_logic;
signal sr_divider_data_7 : std_logic;
signal n8 : std_logic;
signal n3_adj_118 : std_logic;
signal n15 : std_logic;
signal n7 : std_logic;
signal n10 : std_logic;
signal n14 : std_logic;
signal n2_adj_99 : std_logic;
signal n11 : std_logic;
signal \n823_cascade_\ : std_logic;
signal n781 : std_logic;
signal n827 : std_logic;
signal sr_sel_row_c : std_logic;
signal \n169_cascade_\ : std_logic;
signal sr_sel_div_c : std_logic;
signal sr_reset_c : std_logic;
signal \n330_cascade_\ : std_logic;
signal shifted_data_14 : std_logic;
signal shifted_data_15 : std_logic;
signal shifted_data_11 : std_logic;
signal shifted_data_12 : std_logic;
signal shifted_data_13 : std_logic;
signal shifted_data_8 : std_logic;
signal shifted_data_9 : std_logic;
signal shifted_data_10 : std_logic;
signal shifted_data_5 : std_logic;
signal shifted_data_6 : std_logic;
signal shifted_data_7 : std_logic;
signal \bfn_5_7_0_\ : std_logic;
signal \row_counter.n743\ : std_logic;
signal \row_counter.n744\ : std_logic;
signal \row_counter.n745\ : std_logic;
signal \row_counter.n746\ : std_logic;
signal \row_counter.n747\ : std_logic;
signal \row_counter.n748\ : std_logic;
signal \row_counter.n749\ : std_logic;
signal \row_counter.n750\ : std_logic;
signal \bfn_5_8_0_\ : std_logic;
signal \row_counter.n751\ : std_logic;
signal \row_counter.n752\ : std_logic;
signal \row_counter.n753\ : std_logic;
signal \row_counter.n754\ : std_logic;
signal \row_counter.n755\ : std_logic;
signal \row_counter.n756\ : std_logic;
signal \row_counter.n757\ : std_logic;
signal en_rowpack_c : std_logic;
signal n189 : std_logic;
signal sr_data_c : std_logic;
signal shifted_data_0 : std_logic;
signal shifted_data_1 : std_logic;
signal shifted_data_2 : std_logic;
signal n330 : std_logic;
signal n169 : std_logic;
signal shifted_data_3 : std_logic;
signal shifted_data_4 : std_logic;
signal shifted_data_0_adj_115 : std_logic;
signal shifted_data_1_adj_114 : std_logic;
signal \row_counter.internal_count_0\ : std_logic;
signal sr_row_data_0 : std_logic;
signal \bfn_6_7_0_\ : std_logic;
signal \row_counter.internal_count_1\ : std_logic;
signal sr_row_data_1 : std_logic;
signal \row_counter.n696\ : std_logic;
signal \row_counter.internal_count_2\ : std_logic;
signal \row_counter.n697\ : std_logic;
signal \row_counter.internal_count_3\ : std_logic;
signal \row_counter.n698\ : std_logic;
signal \row_counter.internal_count_4\ : std_logic;
signal sr_row_data_4 : std_logic;
signal \row_counter.n699\ : std_logic;
signal \row_counter.internal_count_5\ : std_logic;
signal \row_counter.n700\ : std_logic;
signal \row_counter.internal_count_6\ : std_logic;
signal \row_counter.n701\ : std_logic;
signal \row_counter.internal_count_7\ : std_logic;
signal sr_row_data_7 : std_logic;
signal \row_counter.n702\ : std_logic;
signal \row_counter.n703\ : std_logic;
signal \row_counter.internal_count_8\ : std_logic;
signal \bfn_6_8_0_\ : std_logic;
signal \row_counter.internal_count_9\ : std_logic;
signal \row_counter.n704\ : std_logic;
signal \row_counter.internal_count_10\ : std_logic;
signal \row_counter.n705\ : std_logic;
signal \row_counter.internal_count_11\ : std_logic;
signal \row_counter.n706\ : std_logic;
signal \row_counter.internal_count_12\ : std_logic;
signal \row_counter.n707\ : std_logic;
signal \row_counter.internal_count_13\ : std_logic;
signal \row_counter.n708\ : std_logic;
signal \row_counter.internal_count_14\ : std_logic;
signal \row_counter.n709\ : std_logic;
signal \row_counter.internal_count_15\ : std_logic;
signal \row_counter.n710\ : std_logic;
signal \row_counter.n711\ : std_logic;
signal \row_counter.n13\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \bfn_6_9_0_\ : std_logic;
signal sr_row_data_8 : std_logic;
signal sr_row_data_6 : std_logic;
signal sr_row_data_9 : std_logic;
signal n4 : std_logic;
signal n5 : std_logic;
signal n1 : std_logic;
signal n9_adj_123 : std_logic;
signal \n811_cascade_\ : std_logic;
signal n6 : std_logic;
signal n12_adj_126 : std_logic;
signal n16_adj_129 : std_logic;
signal \n831_cascade_\ : std_logic;
signal n775 : std_logic;
signal reset_signal : std_logic;
signal \n835_cascade_\ : std_logic;
signal row_complete : std_logic;
signal divided_pulse_c : std_logic;
signal sr_row_data_14 : std_logic;
signal sr_row_data_11 : std_logic;
signal sr_row_data_15 : std_logic;
signal sr_row_data_13 : std_logic;
signal shifted_data_15_adj_100 : std_logic;
signal shifted_data_14_adj_101 : std_logic;
signal sr_row_data_10 : std_logic;
signal shifted_data_2_adj_113 : std_logic;
signal sr_row_data_2 : std_logic;
signal n8_adj_122 : std_logic;
signal n3 : std_logic;
signal shifted_data_4_adj_111 : std_logic;
signal n15_adj_128 : std_logic;
signal n7_adj_121 : std_logic;
signal n10_adj_124 : std_logic;
signal n14_adj_127 : std_logic;
signal n2 : std_logic;
signal n11_adj_125 : std_logic;
signal \n793_cascade_\ : std_logic;
signal n803 : std_logic;
signal n829 : std_logic;
signal shifted_data_6_adj_109 : std_logic;
signal shifted_data_7_adj_108 : std_logic;
signal shifted_data_8_adj_107 : std_logic;
signal sr_row_data_12 : std_logic;
signal shifted_data_13_adj_102 : std_logic;
signal shifted_data_11_adj_104 : std_logic;
signal shifted_data_12_adj_103 : std_logic;
signal n345 : std_logic;
signal n171 : std_logic;
signal shifted_data_9_adj_106 : std_logic;
signal shifted_data_10_adj_105 : std_logic;
signal sr_clk_c : std_logic;
signal shifted_data_5_adj_110 : std_logic;
signal sr_row_data_5 : std_logic;
signal en_internals_c : std_logic;
signal shifted_data_3_adj_112 : std_logic;
signal sr_row_data_3 : std_logic;
signal \_gnd_net_\ : std_logic;

signal sr_clk_wire : std_logic;
signal laser_pulse_wire : std_logic;
signal en_internals_wire : std_logic;
signal sr_reset_wire : std_logic;
signal sr_data_wire : std_logic;
signal divide_enable_wire : std_logic;
signal sr_sel_div_wire : std_logic;
signal constant_v_wire : std_logic;
signal divided_pulse_wire : std_logic;
signal en_rowpack_wire : std_logic;
signal sr_sel_row_wire : std_logic;
signal row_completed_wire : std_logic;

begin
    sr_clk_wire <= sr_clk;
    laser_pulse_wire <= laser_pulse;
    en_internals_wire <= en_internals;
    sr_reset_wire <= sr_reset;
    sr_data_wire <= sr_data;
    divide_enable_wire <= divide_enable;
    sr_sel_div_wire <= sr_sel_div;
    constant_v_wire <= constant_v;
    divided_pulse <= divided_pulse_wire;
    en_rowpack_wire <= en_rowpack;
    sr_sel_row_wire <= sr_sel_row;
    row_completed <= row_completed_wire;

    \sr_clk_pad_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__5168\,
            GLOBALBUFFEROUTPUT => sr_clk_c
        );

    \sr_clk_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5170\,
            DIN => \N__5169\,
            DOUT => \N__5168\,
            PACKAGEPIN => sr_clk_wire
        );

    \sr_clk_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5170\,
            PADOUT => \N__5169\,
            PADIN => \N__5168\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \laser_pulse_pad_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__5158\,
            GLOBALBUFFEROUTPUT => laser_pulse_c
        );

    \laser_pulse_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5160\,
            DIN => \N__5159\,
            DOUT => \N__5158\,
            PACKAGEPIN => laser_pulse_wire
        );

    \laser_pulse_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5160\,
            PADOUT => \N__5159\,
            PADIN => \N__5158\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \en_internals_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5149\,
            DIN => \N__5148\,
            DOUT => \N__5147\,
            PACKAGEPIN => en_internals_wire
        );

    \en_internals_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5149\,
            PADOUT => \N__5148\,
            PADIN => \N__5147\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => en_internals_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \sr_reset_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5140\,
            DIN => \N__5139\,
            DOUT => \N__5138\,
            PACKAGEPIN => sr_reset_wire
        );

    \sr_reset_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5140\,
            PADOUT => \N__5139\,
            PADIN => \N__5138\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => sr_reset_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \sr_data_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5131\,
            DIN => \N__5130\,
            DOUT => \N__5129\,
            PACKAGEPIN => sr_data_wire
        );

    \sr_data_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5131\,
            PADOUT => \N__5130\,
            PADIN => \N__5129\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => sr_data_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \divide_enable_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5122\,
            DIN => \N__5121\,
            DOUT => \N__5120\,
            PACKAGEPIN => divide_enable_wire
        );

    \divide_enable_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5122\,
            PADOUT => \N__5121\,
            PADIN => \N__5120\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => divide_enable_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \sr_sel_div_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5113\,
            DIN => \N__5112\,
            DOUT => \N__5111\,
            PACKAGEPIN => sr_sel_div_wire
        );

    \sr_sel_div_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5113\,
            PADOUT => \N__5112\,
            PADIN => \N__5111\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => sr_sel_div_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \constant_v_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5104\,
            DIN => \N__5103\,
            DOUT => \N__5102\,
            PACKAGEPIN => constant_v_wire
        );

    \constant_v_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5104\,
            PADOUT => \N__5103\,
            PADIN => \N__5102\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => constant_v_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \divided_pulse_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5095\,
            DIN => \N__5094\,
            DOUT => \N__5093\,
            PACKAGEPIN => divided_pulse_wire
        );

    \divided_pulse_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5095\,
            PADOUT => \N__5094\,
            PADIN => \N__5093\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3789\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \en_rowpack_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5086\,
            DIN => \N__5085\,
            DOUT => \N__5084\,
            PACKAGEPIN => en_rowpack_wire
        );

    \en_rowpack_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5086\,
            PADOUT => \N__5085\,
            PADIN => \N__5084\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => en_rowpack_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \sr_sel_row_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5077\,
            DIN => \N__5076\,
            DOUT => \N__5075\,
            PACKAGEPIN => sr_sel_row_wire
        );

    \sr_sel_row_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5077\,
            PADOUT => \N__5076\,
            PADIN => \N__5075\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => sr_sel_row_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \row_completed_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5068\,
            DIN => \N__5067\,
            DOUT => \N__5066\,
            PACKAGEPIN => row_completed_wire
        );

    \row_completed_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5068\,
            PADOUT => \N__5067\,
            PADIN => \N__5066\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1164\ : InMux
    port map (
            O => \N__5049\,
            I => \N__5044\
        );

    \I__1163\ : InMux
    port map (
            O => \N__5048\,
            I => \N__5039\
        );

    \I__1162\ : InMux
    port map (
            O => \N__5047\,
            I => \N__5039\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__5044\,
            I => shifted_data_8_adj_107
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__5039\,
            I => shifted_data_8_adj_107
        );

    \I__1159\ : InMux
    port map (
            O => \N__5034\,
            I => \N__5031\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__5031\,
            I => \N__5028\
        );

    \I__1157\ : Odrv4
    port map (
            O => \N__5028\,
            I => sr_row_data_12
        );

    \I__1156\ : CascadeMux
    port map (
            O => \N__5025\,
            I => \N__5020\
        );

    \I__1155\ : InMux
    port map (
            O => \N__5024\,
            I => \N__5015\
        );

    \I__1154\ : InMux
    port map (
            O => \N__5023\,
            I => \N__5015\
        );

    \I__1153\ : InMux
    port map (
            O => \N__5020\,
            I => \N__5012\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__5015\,
            I => shifted_data_13_adj_102
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__5012\,
            I => shifted_data_13_adj_102
        );

    \I__1150\ : CascadeMux
    port map (
            O => \N__5007\,
            I => \N__5004\
        );

    \I__1149\ : InMux
    port map (
            O => \N__5004\,
            I => \N__4999\
        );

    \I__1148\ : InMux
    port map (
            O => \N__5003\,
            I => \N__4994\
        );

    \I__1147\ : InMux
    port map (
            O => \N__5002\,
            I => \N__4994\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__4999\,
            I => shifted_data_11_adj_104
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__4994\,
            I => shifted_data_11_adj_104
        );

    \I__1144\ : InMux
    port map (
            O => \N__4989\,
            I => \N__4980\
        );

    \I__1143\ : InMux
    port map (
            O => \N__4988\,
            I => \N__4980\
        );

    \I__1142\ : InMux
    port map (
            O => \N__4987\,
            I => \N__4980\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__4980\,
            I => shifted_data_12_adj_103
        );

    \I__1140\ : CascadeMux
    port map (
            O => \N__4977\,
            I => \N__4972\
        );

    \I__1139\ : InMux
    port map (
            O => \N__4976\,
            I => \N__4958\
        );

    \I__1138\ : InMux
    port map (
            O => \N__4975\,
            I => \N__4951\
        );

    \I__1137\ : InMux
    port map (
            O => \N__4972\,
            I => \N__4951\
        );

    \I__1136\ : InMux
    port map (
            O => \N__4971\,
            I => \N__4951\
        );

    \I__1135\ : InMux
    port map (
            O => \N__4970\,
            I => \N__4948\
        );

    \I__1134\ : InMux
    port map (
            O => \N__4969\,
            I => \N__4941\
        );

    \I__1133\ : InMux
    port map (
            O => \N__4968\,
            I => \N__4941\
        );

    \I__1132\ : InMux
    port map (
            O => \N__4967\,
            I => \N__4941\
        );

    \I__1131\ : InMux
    port map (
            O => \N__4966\,
            I => \N__4936\
        );

    \I__1130\ : InMux
    port map (
            O => \N__4965\,
            I => \N__4936\
        );

    \I__1129\ : InMux
    port map (
            O => \N__4964\,
            I => \N__4933\
        );

    \I__1128\ : InMux
    port map (
            O => \N__4963\,
            I => \N__4926\
        );

    \I__1127\ : InMux
    port map (
            O => \N__4962\,
            I => \N__4926\
        );

    \I__1126\ : InMux
    port map (
            O => \N__4961\,
            I => \N__4926\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__4958\,
            I => \N__4917\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__4951\,
            I => \N__4917\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__4948\,
            I => \N__4917\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__4941\,
            I => \N__4914\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__4936\,
            I => \N__4909\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__4933\,
            I => \N__4909\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__4926\,
            I => \N__4906\
        );

    \I__1118\ : InMux
    port map (
            O => \N__4925\,
            I => \N__4901\
        );

    \I__1117\ : InMux
    port map (
            O => \N__4924\,
            I => \N__4901\
        );

    \I__1116\ : Span4Mux_v
    port map (
            O => \N__4917\,
            I => \N__4896\
        );

    \I__1115\ : Span4Mux_v
    port map (
            O => \N__4914\,
            I => \N__4896\
        );

    \I__1114\ : Span4Mux_v
    port map (
            O => \N__4909\,
            I => \N__4891\
        );

    \I__1113\ : Span4Mux_v
    port map (
            O => \N__4906\,
            I => \N__4891\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__4901\,
            I => \N__4888\
        );

    \I__1111\ : Odrv4
    port map (
            O => \N__4896\,
            I => n345
        );

    \I__1110\ : Odrv4
    port map (
            O => \N__4891\,
            I => n345
        );

    \I__1109\ : Odrv12
    port map (
            O => \N__4888\,
            I => n345
        );

    \I__1108\ : CascadeMux
    port map (
            O => \N__4881\,
            I => \N__4873\
        );

    \I__1107\ : CascadeMux
    port map (
            O => \N__4880\,
            I => \N__4868\
        );

    \I__1106\ : CascadeMux
    port map (
            O => \N__4879\,
            I => \N__4865\
        );

    \I__1105\ : CascadeMux
    port map (
            O => \N__4878\,
            I => \N__4859\
        );

    \I__1104\ : CascadeMux
    port map (
            O => \N__4877\,
            I => \N__4856\
        );

    \I__1103\ : CascadeMux
    port map (
            O => \N__4876\,
            I => \N__4853\
        );

    \I__1102\ : InMux
    port map (
            O => \N__4873\,
            I => \N__4846\
        );

    \I__1101\ : InMux
    port map (
            O => \N__4872\,
            I => \N__4846\
        );

    \I__1100\ : InMux
    port map (
            O => \N__4871\,
            I => \N__4846\
        );

    \I__1099\ : InMux
    port map (
            O => \N__4868\,
            I => \N__4841\
        );

    \I__1098\ : InMux
    port map (
            O => \N__4865\,
            I => \N__4841\
        );

    \I__1097\ : CascadeMux
    port map (
            O => \N__4864\,
            I => \N__4836\
        );

    \I__1096\ : CascadeMux
    port map (
            O => \N__4863\,
            I => \N__4832\
        );

    \I__1095\ : CascadeMux
    port map (
            O => \N__4862\,
            I => \N__4829\
        );

    \I__1094\ : InMux
    port map (
            O => \N__4859\,
            I => \N__4825\
        );

    \I__1093\ : InMux
    port map (
            O => \N__4856\,
            I => \N__4822\
        );

    \I__1092\ : InMux
    port map (
            O => \N__4853\,
            I => \N__4819\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__4846\,
            I => \N__4814\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__4841\,
            I => \N__4814\
        );

    \I__1089\ : InMux
    port map (
            O => \N__4840\,
            I => \N__4809\
        );

    \I__1088\ : InMux
    port map (
            O => \N__4839\,
            I => \N__4809\
        );

    \I__1087\ : InMux
    port map (
            O => \N__4836\,
            I => \N__4806\
        );

    \I__1086\ : InMux
    port map (
            O => \N__4835\,
            I => \N__4799\
        );

    \I__1085\ : InMux
    port map (
            O => \N__4832\,
            I => \N__4799\
        );

    \I__1084\ : InMux
    port map (
            O => \N__4829\,
            I => \N__4799\
        );

    \I__1083\ : CascadeMux
    port map (
            O => \N__4828\,
            I => \N__4795\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__4825\,
            I => \N__4792\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__4822\,
            I => \N__4787\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__4819\,
            I => \N__4787\
        );

    \I__1079\ : Span4Mux_v
    port map (
            O => \N__4814\,
            I => \N__4778\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__4809\,
            I => \N__4778\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__4806\,
            I => \N__4778\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__4799\,
            I => \N__4778\
        );

    \I__1075\ : InMux
    port map (
            O => \N__4798\,
            I => \N__4773\
        );

    \I__1074\ : InMux
    port map (
            O => \N__4795\,
            I => \N__4773\
        );

    \I__1073\ : Span4Mux_v
    port map (
            O => \N__4792\,
            I => \N__4770\
        );

    \I__1072\ : Span4Mux_v
    port map (
            O => \N__4787\,
            I => \N__4765\
        );

    \I__1071\ : Span4Mux_v
    port map (
            O => \N__4778\,
            I => \N__4765\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__4773\,
            I => \N__4762\
        );

    \I__1069\ : Odrv4
    port map (
            O => \N__4770\,
            I => n171
        );

    \I__1068\ : Odrv4
    port map (
            O => \N__4765\,
            I => n171
        );

    \I__1067\ : Odrv12
    port map (
            O => \N__4762\,
            I => n171
        );

    \I__1066\ : CascadeMux
    port map (
            O => \N__4755\,
            I => \N__4750\
        );

    \I__1065\ : InMux
    port map (
            O => \N__4754\,
            I => \N__4747\
        );

    \I__1064\ : InMux
    port map (
            O => \N__4753\,
            I => \N__4744\
        );

    \I__1063\ : InMux
    port map (
            O => \N__4750\,
            I => \N__4741\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__4747\,
            I => shifted_data_9_adj_106
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__4744\,
            I => shifted_data_9_adj_106
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__4741\,
            I => shifted_data_9_adj_106
        );

    \I__1059\ : InMux
    port map (
            O => \N__4734\,
            I => \N__4727\
        );

    \I__1058\ : InMux
    port map (
            O => \N__4733\,
            I => \N__4727\
        );

    \I__1057\ : InMux
    port map (
            O => \N__4732\,
            I => \N__4724\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__4727\,
            I => shifted_data_10_adj_105
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__4724\,
            I => shifted_data_10_adj_105
        );

    \I__1054\ : ClkMux
    port map (
            O => \N__4719\,
            I => \N__4683\
        );

    \I__1053\ : ClkMux
    port map (
            O => \N__4718\,
            I => \N__4683\
        );

    \I__1052\ : ClkMux
    port map (
            O => \N__4717\,
            I => \N__4683\
        );

    \I__1051\ : ClkMux
    port map (
            O => \N__4716\,
            I => \N__4683\
        );

    \I__1050\ : ClkMux
    port map (
            O => \N__4715\,
            I => \N__4683\
        );

    \I__1049\ : ClkMux
    port map (
            O => \N__4714\,
            I => \N__4683\
        );

    \I__1048\ : ClkMux
    port map (
            O => \N__4713\,
            I => \N__4683\
        );

    \I__1047\ : ClkMux
    port map (
            O => \N__4712\,
            I => \N__4683\
        );

    \I__1046\ : ClkMux
    port map (
            O => \N__4711\,
            I => \N__4683\
        );

    \I__1045\ : ClkMux
    port map (
            O => \N__4710\,
            I => \N__4683\
        );

    \I__1044\ : ClkMux
    port map (
            O => \N__4709\,
            I => \N__4683\
        );

    \I__1043\ : ClkMux
    port map (
            O => \N__4708\,
            I => \N__4683\
        );

    \I__1042\ : GlobalMux
    port map (
            O => \N__4683\,
            I => \N__4680\
        );

    \I__1041\ : gio2CtrlBuf
    port map (
            O => \N__4680\,
            I => sr_clk_c
        );

    \I__1040\ : InMux
    port map (
            O => \N__4677\,
            I => \N__4672\
        );

    \I__1039\ : InMux
    port map (
            O => \N__4676\,
            I => \N__4667\
        );

    \I__1038\ : InMux
    port map (
            O => \N__4675\,
            I => \N__4667\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__4672\,
            I => shifted_data_5_adj_110
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__4667\,
            I => shifted_data_5_adj_110
        );

    \I__1035\ : CascadeMux
    port map (
            O => \N__4662\,
            I => \N__4659\
        );

    \I__1034\ : InMux
    port map (
            O => \N__4659\,
            I => \N__4656\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__4656\,
            I => \N__4653\
        );

    \I__1032\ : Odrv4
    port map (
            O => \N__4653\,
            I => sr_row_data_5
        );

    \I__1031\ : InMux
    port map (
            O => \N__4650\,
            I => \N__4642\
        );

    \I__1030\ : InMux
    port map (
            O => \N__4649\,
            I => \N__4639\
        );

    \I__1029\ : InMux
    port map (
            O => \N__4648\,
            I => \N__4632\
        );

    \I__1028\ : InMux
    port map (
            O => \N__4647\,
            I => \N__4632\
        );

    \I__1027\ : InMux
    port map (
            O => \N__4646\,
            I => \N__4632\
        );

    \I__1026\ : InMux
    port map (
            O => \N__4645\,
            I => \N__4624\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__4642\,
            I => \N__4612\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__4639\,
            I => \N__4612\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__4632\,
            I => \N__4612\
        );

    \I__1022\ : InMux
    port map (
            O => \N__4631\,
            I => \N__4601\
        );

    \I__1021\ : InMux
    port map (
            O => \N__4630\,
            I => \N__4601\
        );

    \I__1020\ : InMux
    port map (
            O => \N__4629\,
            I => \N__4601\
        );

    \I__1019\ : InMux
    port map (
            O => \N__4628\,
            I => \N__4601\
        );

    \I__1018\ : InMux
    port map (
            O => \N__4627\,
            I => \N__4601\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__4624\,
            I => \N__4598\
        );

    \I__1016\ : InMux
    port map (
            O => \N__4623\,
            I => \N__4593\
        );

    \I__1015\ : InMux
    port map (
            O => \N__4622\,
            I => \N__4593\
        );

    \I__1014\ : InMux
    port map (
            O => \N__4621\,
            I => \N__4578\
        );

    \I__1013\ : InMux
    port map (
            O => \N__4620\,
            I => \N__4578\
        );

    \I__1012\ : InMux
    port map (
            O => \N__4619\,
            I => \N__4578\
        );

    \I__1011\ : Span4Mux_v
    port map (
            O => \N__4612\,
            I => \N__4573\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__4601\,
            I => \N__4573\
        );

    \I__1009\ : Span4Mux_h
    port map (
            O => \N__4598\,
            I => \N__4568\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__4593\,
            I => \N__4568\
        );

    \I__1007\ : InMux
    port map (
            O => \N__4592\,
            I => \N__4551\
        );

    \I__1006\ : InMux
    port map (
            O => \N__4591\,
            I => \N__4551\
        );

    \I__1005\ : InMux
    port map (
            O => \N__4590\,
            I => \N__4551\
        );

    \I__1004\ : InMux
    port map (
            O => \N__4589\,
            I => \N__4551\
        );

    \I__1003\ : InMux
    port map (
            O => \N__4588\,
            I => \N__4551\
        );

    \I__1002\ : InMux
    port map (
            O => \N__4587\,
            I => \N__4551\
        );

    \I__1001\ : InMux
    port map (
            O => \N__4586\,
            I => \N__4551\
        );

    \I__1000\ : InMux
    port map (
            O => \N__4585\,
            I => \N__4551\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__4578\,
            I => \N__4540\
        );

    \I__998\ : Span4Mux_h
    port map (
            O => \N__4573\,
            I => \N__4533\
        );

    \I__997\ : Span4Mux_v
    port map (
            O => \N__4568\,
            I => \N__4533\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__4551\,
            I => \N__4533\
        );

    \I__995\ : InMux
    port map (
            O => \N__4550\,
            I => \N__4520\
        );

    \I__994\ : InMux
    port map (
            O => \N__4549\,
            I => \N__4520\
        );

    \I__993\ : InMux
    port map (
            O => \N__4548\,
            I => \N__4520\
        );

    \I__992\ : InMux
    port map (
            O => \N__4547\,
            I => \N__4520\
        );

    \I__991\ : InMux
    port map (
            O => \N__4546\,
            I => \N__4520\
        );

    \I__990\ : InMux
    port map (
            O => \N__4545\,
            I => \N__4520\
        );

    \I__989\ : InMux
    port map (
            O => \N__4544\,
            I => \N__4515\
        );

    \I__988\ : InMux
    port map (
            O => \N__4543\,
            I => \N__4515\
        );

    \I__987\ : Span4Mux_v
    port map (
            O => \N__4540\,
            I => \N__4512\
        );

    \I__986\ : Span4Mux_h
    port map (
            O => \N__4533\,
            I => \N__4507\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__4520\,
            I => \N__4507\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__4515\,
            I => \N__4504\
        );

    \I__983\ : Span4Mux_v
    port map (
            O => \N__4512\,
            I => \N__4501\
        );

    \I__982\ : Span4Mux_v
    port map (
            O => \N__4507\,
            I => \N__4498\
        );

    \I__981\ : Span12Mux_v
    port map (
            O => \N__4504\,
            I => \N__4491\
        );

    \I__980\ : Sp12to4
    port map (
            O => \N__4501\,
            I => \N__4491\
        );

    \I__979\ : Sp12to4
    port map (
            O => \N__4498\,
            I => \N__4491\
        );

    \I__978\ : Odrv12
    port map (
            O => \N__4491\,
            I => en_internals_c
        );

    \I__977\ : CascadeMux
    port map (
            O => \N__4488\,
            I => \N__4485\
        );

    \I__976\ : InMux
    port map (
            O => \N__4485\,
            I => \N__4481\
        );

    \I__975\ : InMux
    port map (
            O => \N__4484\,
            I => \N__4477\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__4481\,
            I => \N__4474\
        );

    \I__973\ : InMux
    port map (
            O => \N__4480\,
            I => \N__4471\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__4477\,
            I => shifted_data_3_adj_112
        );

    \I__971\ : Odrv4
    port map (
            O => \N__4474\,
            I => shifted_data_3_adj_112
        );

    \I__970\ : LocalMux
    port map (
            O => \N__4471\,
            I => shifted_data_3_adj_112
        );

    \I__969\ : CascadeMux
    port map (
            O => \N__4464\,
            I => \N__4461\
        );

    \I__968\ : InMux
    port map (
            O => \N__4461\,
            I => \N__4458\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__4458\,
            I => \N__4455\
        );

    \I__966\ : Odrv4
    port map (
            O => \N__4455\,
            I => sr_row_data_3
        );

    \I__965\ : InMux
    port map (
            O => \N__4452\,
            I => \N__4447\
        );

    \I__964\ : InMux
    port map (
            O => \N__4451\,
            I => \N__4444\
        );

    \I__963\ : InMux
    port map (
            O => \N__4450\,
            I => \N__4441\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__4447\,
            I => shifted_data_2_adj_113
        );

    \I__961\ : LocalMux
    port map (
            O => \N__4444\,
            I => shifted_data_2_adj_113
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4441\,
            I => shifted_data_2_adj_113
        );

    \I__959\ : InMux
    port map (
            O => \N__4434\,
            I => \N__4431\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__4431\,
            I => sr_row_data_2
        );

    \I__957\ : InMux
    port map (
            O => \N__4428\,
            I => \N__4425\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__4425\,
            I => n8_adj_122
        );

    \I__955\ : InMux
    port map (
            O => \N__4422\,
            I => \N__4419\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__4419\,
            I => n3
        );

    \I__953\ : InMux
    port map (
            O => \N__4416\,
            I => \N__4413\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__4413\,
            I => \N__4410\
        );

    \I__951\ : Span4Mux_v
    port map (
            O => \N__4410\,
            I => \N__4405\
        );

    \I__950\ : InMux
    port map (
            O => \N__4409\,
            I => \N__4400\
        );

    \I__949\ : InMux
    port map (
            O => \N__4408\,
            I => \N__4400\
        );

    \I__948\ : Odrv4
    port map (
            O => \N__4405\,
            I => shifted_data_4_adj_111
        );

    \I__947\ : LocalMux
    port map (
            O => \N__4400\,
            I => shifted_data_4_adj_111
        );

    \I__946\ : InMux
    port map (
            O => \N__4395\,
            I => \N__4392\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__4392\,
            I => n15_adj_128
        );

    \I__944\ : InMux
    port map (
            O => \N__4389\,
            I => \N__4386\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__4386\,
            I => n7_adj_121
        );

    \I__942\ : CascadeMux
    port map (
            O => \N__4383\,
            I => \N__4380\
        );

    \I__941\ : InMux
    port map (
            O => \N__4380\,
            I => \N__4377\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__4377\,
            I => n10_adj_124
        );

    \I__939\ : InMux
    port map (
            O => \N__4374\,
            I => \N__4371\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__4371\,
            I => n14_adj_127
        );

    \I__937\ : InMux
    port map (
            O => \N__4368\,
            I => \N__4365\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__4365\,
            I => n2
        );

    \I__935\ : InMux
    port map (
            O => \N__4362\,
            I => \N__4359\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__4359\,
            I => n11_adj_125
        );

    \I__933\ : CascadeMux
    port map (
            O => \N__4356\,
            I => \n793_cascade_\
        );

    \I__932\ : InMux
    port map (
            O => \N__4353\,
            I => \N__4350\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__4350\,
            I => n803
        );

    \I__930\ : InMux
    port map (
            O => \N__4347\,
            I => \N__4344\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__4344\,
            I => n829
        );

    \I__928\ : InMux
    port map (
            O => \N__4341\,
            I => \N__4338\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__4338\,
            I => \N__4333\
        );

    \I__926\ : InMux
    port map (
            O => \N__4337\,
            I => \N__4330\
        );

    \I__925\ : InMux
    port map (
            O => \N__4336\,
            I => \N__4327\
        );

    \I__924\ : Odrv4
    port map (
            O => \N__4333\,
            I => shifted_data_6_adj_109
        );

    \I__923\ : LocalMux
    port map (
            O => \N__4330\,
            I => shifted_data_6_adj_109
        );

    \I__922\ : LocalMux
    port map (
            O => \N__4327\,
            I => shifted_data_6_adj_109
        );

    \I__921\ : InMux
    port map (
            O => \N__4320\,
            I => \N__4317\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__4317\,
            I => \N__4314\
        );

    \I__919\ : Span4Mux_v
    port map (
            O => \N__4314\,
            I => \N__4309\
        );

    \I__918\ : InMux
    port map (
            O => \N__4313\,
            I => \N__4306\
        );

    \I__917\ : InMux
    port map (
            O => \N__4312\,
            I => \N__4303\
        );

    \I__916\ : Odrv4
    port map (
            O => \N__4309\,
            I => shifted_data_7_adj_108
        );

    \I__915\ : LocalMux
    port map (
            O => \N__4306\,
            I => shifted_data_7_adj_108
        );

    \I__914\ : LocalMux
    port map (
            O => \N__4303\,
            I => shifted_data_7_adj_108
        );

    \I__913\ : InMux
    port map (
            O => \N__4296\,
            I => \N__4293\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__4293\,
            I => \N__4290\
        );

    \I__911\ : Odrv4
    port map (
            O => \N__4290\,
            I => sr_row_data_14
        );

    \I__910\ : InMux
    port map (
            O => \N__4287\,
            I => \N__4284\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__4284\,
            I => \N__4281\
        );

    \I__908\ : Odrv4
    port map (
            O => \N__4281\,
            I => sr_row_data_11
        );

    \I__907\ : InMux
    port map (
            O => \N__4278\,
            I => \N__4275\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__4275\,
            I => \N__4272\
        );

    \I__905\ : Odrv4
    port map (
            O => \N__4272\,
            I => sr_row_data_15
        );

    \I__904\ : InMux
    port map (
            O => \N__4269\,
            I => \N__4266\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__4266\,
            I => \N__4263\
        );

    \I__902\ : Odrv4
    port map (
            O => \N__4263\,
            I => sr_row_data_13
        );

    \I__901\ : CascadeMux
    port map (
            O => \N__4260\,
            I => \N__4256\
        );

    \I__900\ : InMux
    port map (
            O => \N__4259\,
            I => \N__4251\
        );

    \I__899\ : InMux
    port map (
            O => \N__4256\,
            I => \N__4251\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__4251\,
            I => shifted_data_15_adj_100
        );

    \I__897\ : InMux
    port map (
            O => \N__4248\,
            I => \N__4239\
        );

    \I__896\ : InMux
    port map (
            O => \N__4247\,
            I => \N__4239\
        );

    \I__895\ : InMux
    port map (
            O => \N__4246\,
            I => \N__4239\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__4239\,
            I => shifted_data_14_adj_101
        );

    \I__893\ : InMux
    port map (
            O => \N__4236\,
            I => \N__4233\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__4233\,
            I => \N__4230\
        );

    \I__891\ : Odrv4
    port map (
            O => \N__4230\,
            I => sr_row_data_10
        );

    \I__890\ : InMux
    port map (
            O => \N__4227\,
            I => \N__4224\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__4224\,
            I => \row_counter.n13\
        );

    \I__888\ : CascadeMux
    port map (
            O => \N__4221\,
            I => \N__4209\
        );

    \I__887\ : CascadeMux
    port map (
            O => \N__4220\,
            I => \N__4206\
        );

    \I__886\ : CascadeMux
    port map (
            O => \N__4219\,
            I => \N__4202\
        );

    \I__885\ : CascadeMux
    port map (
            O => \N__4218\,
            I => \N__4198\
        );

    \I__884\ : CascadeMux
    port map (
            O => \N__4217\,
            I => \N__4194\
        );

    \I__883\ : CascadeMux
    port map (
            O => \N__4216\,
            I => \N__4191\
        );

    \I__882\ : CascadeMux
    port map (
            O => \N__4215\,
            I => \N__4186\
        );

    \I__881\ : CascadeMux
    port map (
            O => \N__4214\,
            I => \N__4183\
        );

    \I__880\ : CascadeMux
    port map (
            O => \N__4213\,
            I => \N__4180\
        );

    \I__879\ : CascadeMux
    port map (
            O => \N__4212\,
            I => \N__4177\
        );

    \I__878\ : InMux
    port map (
            O => \N__4209\,
            I => \N__4164\
        );

    \I__877\ : InMux
    port map (
            O => \N__4206\,
            I => \N__4164\
        );

    \I__876\ : InMux
    port map (
            O => \N__4205\,
            I => \N__4164\
        );

    \I__875\ : InMux
    port map (
            O => \N__4202\,
            I => \N__4164\
        );

    \I__874\ : InMux
    port map (
            O => \N__4201\,
            I => \N__4164\
        );

    \I__873\ : InMux
    port map (
            O => \N__4198\,
            I => \N__4164\
        );

    \I__872\ : InMux
    port map (
            O => \N__4197\,
            I => \N__4157\
        );

    \I__871\ : InMux
    port map (
            O => \N__4194\,
            I => \N__4157\
        );

    \I__870\ : InMux
    port map (
            O => \N__4191\,
            I => \N__4157\
        );

    \I__869\ : InMux
    port map (
            O => \N__4190\,
            I => \N__4146\
        );

    \I__868\ : InMux
    port map (
            O => \N__4189\,
            I => \N__4146\
        );

    \I__867\ : InMux
    port map (
            O => \N__4186\,
            I => \N__4146\
        );

    \I__866\ : InMux
    port map (
            O => \N__4183\,
            I => \N__4146\
        );

    \I__865\ : InMux
    port map (
            O => \N__4180\,
            I => \N__4146\
        );

    \I__864\ : InMux
    port map (
            O => \N__4177\,
            I => \N__4140\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__4164\,
            I => \N__4133\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__4157\,
            I => \N__4133\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__4146\,
            I => \N__4133\
        );

    \I__860\ : CascadeMux
    port map (
            O => \N__4145\,
            I => \N__4129\
        );

    \I__859\ : CascadeMux
    port map (
            O => \N__4144\,
            I => \N__4125\
        );

    \I__858\ : CascadeMux
    port map (
            O => \N__4143\,
            I => \N__4121\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__4140\,
            I => \N__4108\
        );

    \I__856\ : Span4Mux_v
    port map (
            O => \N__4133\,
            I => \N__4105\
        );

    \I__855\ : InMux
    port map (
            O => \N__4132\,
            I => \N__4090\
        );

    \I__854\ : InMux
    port map (
            O => \N__4129\,
            I => \N__4090\
        );

    \I__853\ : InMux
    port map (
            O => \N__4128\,
            I => \N__4090\
        );

    \I__852\ : InMux
    port map (
            O => \N__4125\,
            I => \N__4090\
        );

    \I__851\ : InMux
    port map (
            O => \N__4124\,
            I => \N__4090\
        );

    \I__850\ : InMux
    port map (
            O => \N__4121\,
            I => \N__4090\
        );

    \I__849\ : InMux
    port map (
            O => \N__4120\,
            I => \N__4090\
        );

    \I__848\ : InMux
    port map (
            O => \N__4119\,
            I => \N__4087\
        );

    \I__847\ : CascadeMux
    port map (
            O => \N__4118\,
            I => \N__4084\
        );

    \I__846\ : CascadeMux
    port map (
            O => \N__4117\,
            I => \N__4081\
        );

    \I__845\ : CascadeMux
    port map (
            O => \N__4116\,
            I => \N__4078\
        );

    \I__844\ : CascadeMux
    port map (
            O => \N__4115\,
            I => \N__4075\
        );

    \I__843\ : CascadeMux
    port map (
            O => \N__4114\,
            I => \N__4072\
        );

    \I__842\ : CascadeMux
    port map (
            O => \N__4113\,
            I => \N__4069\
        );

    \I__841\ : CascadeMux
    port map (
            O => \N__4112\,
            I => \N__4066\
        );

    \I__840\ : CascadeMux
    port map (
            O => \N__4111\,
            I => \N__4063\
        );

    \I__839\ : Span4Mux_v
    port map (
            O => \N__4108\,
            I => \N__4059\
        );

    \I__838\ : Span4Mux_h
    port map (
            O => \N__4105\,
            I => \N__4054\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__4090\,
            I => \N__4054\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__4087\,
            I => \N__4051\
        );

    \I__835\ : InMux
    port map (
            O => \N__4084\,
            I => \N__4042\
        );

    \I__834\ : InMux
    port map (
            O => \N__4081\,
            I => \N__4042\
        );

    \I__833\ : InMux
    port map (
            O => \N__4078\,
            I => \N__4042\
        );

    \I__832\ : InMux
    port map (
            O => \N__4075\,
            I => \N__4042\
        );

    \I__831\ : InMux
    port map (
            O => \N__4072\,
            I => \N__4033\
        );

    \I__830\ : InMux
    port map (
            O => \N__4069\,
            I => \N__4033\
        );

    \I__829\ : InMux
    port map (
            O => \N__4066\,
            I => \N__4033\
        );

    \I__828\ : InMux
    port map (
            O => \N__4063\,
            I => \N__4033\
        );

    \I__827\ : InMux
    port map (
            O => \N__4062\,
            I => \N__4030\
        );

    \I__826\ : Odrv4
    port map (
            O => \N__4059\,
            I => \CONSTANT_ONE_NET\
        );

    \I__825\ : Odrv4
    port map (
            O => \N__4054\,
            I => \CONSTANT_ONE_NET\
        );

    \I__824\ : Odrv12
    port map (
            O => \N__4051\,
            I => \CONSTANT_ONE_NET\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__4042\,
            I => \CONSTANT_ONE_NET\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__4033\,
            I => \CONSTANT_ONE_NET\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__4030\,
            I => \CONSTANT_ONE_NET\
        );

    \I__820\ : InMux
    port map (
            O => \N__4017\,
            I => \bfn_6_9_0_\
        );

    \I__819\ : InMux
    port map (
            O => \N__4014\,
            I => \N__4011\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__4011\,
            I => sr_row_data_8
        );

    \I__817\ : InMux
    port map (
            O => \N__4008\,
            I => \N__4005\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__4005\,
            I => \N__4002\
        );

    \I__815\ : Odrv4
    port map (
            O => \N__4002\,
            I => sr_row_data_6
        );

    \I__814\ : InMux
    port map (
            O => \N__3999\,
            I => \N__3996\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__3996\,
            I => sr_row_data_9
        );

    \I__812\ : InMux
    port map (
            O => \N__3993\,
            I => \N__3990\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__3990\,
            I => \N__3987\
        );

    \I__810\ : Odrv4
    port map (
            O => \N__3987\,
            I => n4
        );

    \I__809\ : InMux
    port map (
            O => \N__3984\,
            I => \N__3981\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__3981\,
            I => \N__3978\
        );

    \I__807\ : Odrv4
    port map (
            O => \N__3978\,
            I => n5
        );

    \I__806\ : InMux
    port map (
            O => \N__3975\,
            I => \N__3972\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__3972\,
            I => \N__3969\
        );

    \I__804\ : Odrv4
    port map (
            O => \N__3969\,
            I => n1
        );

    \I__803\ : InMux
    port map (
            O => \N__3966\,
            I => \N__3963\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__3963\,
            I => n9_adj_123
        );

    \I__801\ : CascadeMux
    port map (
            O => \N__3960\,
            I => \n811_cascade_\
        );

    \I__800\ : InMux
    port map (
            O => \N__3957\,
            I => \N__3954\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__3954\,
            I => \N__3951\
        );

    \I__798\ : Odrv4
    port map (
            O => \N__3951\,
            I => n6
        );

    \I__797\ : InMux
    port map (
            O => \N__3948\,
            I => \N__3945\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__3945\,
            I => \N__3942\
        );

    \I__795\ : Odrv4
    port map (
            O => \N__3942\,
            I => n12_adj_126
        );

    \I__794\ : InMux
    port map (
            O => \N__3939\,
            I => \N__3936\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__3936\,
            I => n16_adj_129
        );

    \I__792\ : CascadeMux
    port map (
            O => \N__3933\,
            I => \n831_cascade_\
        );

    \I__791\ : InMux
    port map (
            O => \N__3930\,
            I => \N__3927\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__3927\,
            I => n775
        );

    \I__789\ : SRMux
    port map (
            O => \N__3924\,
            I => \N__3920\
        );

    \I__788\ : SRMux
    port map (
            O => \N__3923\,
            I => \N__3916\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__3920\,
            I => \N__3910\
        );

    \I__786\ : SRMux
    port map (
            O => \N__3919\,
            I => \N__3907\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__3916\,
            I => \N__3904\
        );

    \I__784\ : SRMux
    port map (
            O => \N__3915\,
            I => \N__3901\
        );

    \I__783\ : InMux
    port map (
            O => \N__3914\,
            I => \N__3898\
        );

    \I__782\ : InMux
    port map (
            O => \N__3913\,
            I => \N__3895\
        );

    \I__781\ : Span4Mux_h
    port map (
            O => \N__3910\,
            I => \N__3886\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__3907\,
            I => \N__3886\
        );

    \I__779\ : Span4Mux_h
    port map (
            O => \N__3904\,
            I => \N__3881\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__3901\,
            I => \N__3881\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__3898\,
            I => \N__3872\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__3895\,
            I => \N__3872\
        );

    \I__775\ : InMux
    port map (
            O => \N__3894\,
            I => \N__3867\
        );

    \I__774\ : InMux
    port map (
            O => \N__3893\,
            I => \N__3867\
        );

    \I__773\ : InMux
    port map (
            O => \N__3892\,
            I => \N__3862\
        );

    \I__772\ : InMux
    port map (
            O => \N__3891\,
            I => \N__3862\
        );

    \I__771\ : Span4Mux_h
    port map (
            O => \N__3886\,
            I => \N__3859\
        );

    \I__770\ : Span4Mux_h
    port map (
            O => \N__3881\,
            I => \N__3856\
        );

    \I__769\ : InMux
    port map (
            O => \N__3880\,
            I => \N__3851\
        );

    \I__768\ : InMux
    port map (
            O => \N__3879\,
            I => \N__3851\
        );

    \I__767\ : InMux
    port map (
            O => \N__3878\,
            I => \N__3846\
        );

    \I__766\ : InMux
    port map (
            O => \N__3877\,
            I => \N__3846\
        );

    \I__765\ : Odrv12
    port map (
            O => \N__3872\,
            I => reset_signal
        );

    \I__764\ : LocalMux
    port map (
            O => \N__3867\,
            I => reset_signal
        );

    \I__763\ : LocalMux
    port map (
            O => \N__3862\,
            I => reset_signal
        );

    \I__762\ : Odrv4
    port map (
            O => \N__3859\,
            I => reset_signal
        );

    \I__761\ : Odrv4
    port map (
            O => \N__3856\,
            I => reset_signal
        );

    \I__760\ : LocalMux
    port map (
            O => \N__3851\,
            I => reset_signal
        );

    \I__759\ : LocalMux
    port map (
            O => \N__3846\,
            I => reset_signal
        );

    \I__758\ : CascadeMux
    port map (
            O => \N__3831\,
            I => \n835_cascade_\
        );

    \I__757\ : InMux
    port map (
            O => \N__3828\,
            I => \N__3825\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__3825\,
            I => \N__3822\
        );

    \I__755\ : Span4Mux_h
    port map (
            O => \N__3822\,
            I => \N__3817\
        );

    \I__754\ : InMux
    port map (
            O => \N__3821\,
            I => \N__3814\
        );

    \I__753\ : InMux
    port map (
            O => \N__3820\,
            I => \N__3811\
        );

    \I__752\ : Odrv4
    port map (
            O => \N__3817\,
            I => row_complete
        );

    \I__751\ : LocalMux
    port map (
            O => \N__3814\,
            I => row_complete
        );

    \I__750\ : LocalMux
    port map (
            O => \N__3811\,
            I => row_complete
        );

    \I__749\ : ClkMux
    port map (
            O => \N__3804\,
            I => \N__3799\
        );

    \I__748\ : ClkMux
    port map (
            O => \N__3803\,
            I => \N__3796\
        );

    \I__747\ : ClkMux
    port map (
            O => \N__3802\,
            I => \N__3793\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__3799\,
            I => \N__3790\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__3796\,
            I => \N__3786\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__3793\,
            I => \N__3783\
        );

    \I__743\ : Span4Mux_v
    port map (
            O => \N__3790\,
            I => \N__3780\
        );

    \I__742\ : IoInMux
    port map (
            O => \N__3789\,
            I => \N__3777\
        );

    \I__741\ : Span4Mux_h
    port map (
            O => \N__3786\,
            I => \N__3774\
        );

    \I__740\ : Span4Mux_h
    port map (
            O => \N__3783\,
            I => \N__3771\
        );

    \I__739\ : Span4Mux_h
    port map (
            O => \N__3780\,
            I => \N__3768\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__3777\,
            I => \N__3765\
        );

    \I__737\ : Odrv4
    port map (
            O => \N__3774\,
            I => divided_pulse_c
        );

    \I__736\ : Odrv4
    port map (
            O => \N__3771\,
            I => divided_pulse_c
        );

    \I__735\ : Odrv4
    port map (
            O => \N__3768\,
            I => divided_pulse_c
        );

    \I__734\ : Odrv12
    port map (
            O => \N__3765\,
            I => divided_pulse_c
        );

    \I__733\ : InMux
    port map (
            O => \N__3756\,
            I => \N__3752\
        );

    \I__732\ : InMux
    port map (
            O => \N__3755\,
            I => \N__3749\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__3752\,
            I => \row_counter.internal_count_8\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__3749\,
            I => \row_counter.internal_count_8\
        );

    \I__729\ : InMux
    port map (
            O => \N__3744\,
            I => \bfn_6_8_0_\
        );

    \I__728\ : InMux
    port map (
            O => \N__3741\,
            I => \N__3737\
        );

    \I__727\ : InMux
    port map (
            O => \N__3740\,
            I => \N__3734\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__3737\,
            I => \N__3731\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__3734\,
            I => \row_counter.internal_count_9\
        );

    \I__724\ : Odrv4
    port map (
            O => \N__3731\,
            I => \row_counter.internal_count_9\
        );

    \I__723\ : InMux
    port map (
            O => \N__3726\,
            I => \row_counter.n704\
        );

    \I__722\ : InMux
    port map (
            O => \N__3723\,
            I => \N__3719\
        );

    \I__721\ : InMux
    port map (
            O => \N__3722\,
            I => \N__3716\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__3719\,
            I => \row_counter.internal_count_10\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__3716\,
            I => \row_counter.internal_count_10\
        );

    \I__718\ : InMux
    port map (
            O => \N__3711\,
            I => \row_counter.n705\
        );

    \I__717\ : InMux
    port map (
            O => \N__3708\,
            I => \N__3704\
        );

    \I__716\ : InMux
    port map (
            O => \N__3707\,
            I => \N__3701\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__3704\,
            I => \row_counter.internal_count_11\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__3701\,
            I => \row_counter.internal_count_11\
        );

    \I__713\ : InMux
    port map (
            O => \N__3696\,
            I => \row_counter.n706\
        );

    \I__712\ : InMux
    port map (
            O => \N__3693\,
            I => \N__3689\
        );

    \I__711\ : InMux
    port map (
            O => \N__3692\,
            I => \N__3686\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__3689\,
            I => \row_counter.internal_count_12\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__3686\,
            I => \row_counter.internal_count_12\
        );

    \I__708\ : InMux
    port map (
            O => \N__3681\,
            I => \row_counter.n707\
        );

    \I__707\ : InMux
    port map (
            O => \N__3678\,
            I => \N__3674\
        );

    \I__706\ : InMux
    port map (
            O => \N__3677\,
            I => \N__3671\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__3674\,
            I => \row_counter.internal_count_13\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__3671\,
            I => \row_counter.internal_count_13\
        );

    \I__703\ : InMux
    port map (
            O => \N__3666\,
            I => \row_counter.n708\
        );

    \I__702\ : InMux
    port map (
            O => \N__3663\,
            I => \N__3659\
        );

    \I__701\ : InMux
    port map (
            O => \N__3662\,
            I => \N__3656\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__3659\,
            I => \row_counter.internal_count_14\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__3656\,
            I => \row_counter.internal_count_14\
        );

    \I__698\ : InMux
    port map (
            O => \N__3651\,
            I => \row_counter.n709\
        );

    \I__697\ : InMux
    port map (
            O => \N__3648\,
            I => \N__3644\
        );

    \I__696\ : InMux
    port map (
            O => \N__3647\,
            I => \N__3641\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__3644\,
            I => \row_counter.internal_count_15\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__3641\,
            I => \row_counter.internal_count_15\
        );

    \I__693\ : InMux
    port map (
            O => \N__3636\,
            I => \row_counter.n710\
        );

    \I__692\ : InMux
    port map (
            O => \N__3633\,
            I => \N__3624\
        );

    \I__691\ : InMux
    port map (
            O => \N__3632\,
            I => \N__3624\
        );

    \I__690\ : InMux
    port map (
            O => \N__3631\,
            I => \N__3624\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__3624\,
            I => shifted_data_1_adj_114
        );

    \I__688\ : InMux
    port map (
            O => \N__3621\,
            I => \N__3617\
        );

    \I__687\ : InMux
    port map (
            O => \N__3620\,
            I => \N__3614\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__3617\,
            I => \row_counter.internal_count_0\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__3614\,
            I => \row_counter.internal_count_0\
        );

    \I__684\ : InMux
    port map (
            O => \N__3609\,
            I => \N__3606\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__3606\,
            I => \N__3603\
        );

    \I__682\ : Odrv4
    port map (
            O => \N__3603\,
            I => sr_row_data_0
        );

    \I__681\ : InMux
    port map (
            O => \N__3600\,
            I => \bfn_6_7_0_\
        );

    \I__680\ : InMux
    port map (
            O => \N__3597\,
            I => \N__3593\
        );

    \I__679\ : InMux
    port map (
            O => \N__3596\,
            I => \N__3590\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__3593\,
            I => \row_counter.internal_count_1\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__3590\,
            I => \row_counter.internal_count_1\
        );

    \I__676\ : CascadeMux
    port map (
            O => \N__3585\,
            I => \N__3582\
        );

    \I__675\ : InMux
    port map (
            O => \N__3582\,
            I => \N__3579\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__3579\,
            I => sr_row_data_1
        );

    \I__673\ : InMux
    port map (
            O => \N__3576\,
            I => \row_counter.n696\
        );

    \I__672\ : InMux
    port map (
            O => \N__3573\,
            I => \N__3569\
        );

    \I__671\ : InMux
    port map (
            O => \N__3572\,
            I => \N__3566\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__3569\,
            I => \N__3561\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__3566\,
            I => \N__3561\
        );

    \I__668\ : Odrv4
    port map (
            O => \N__3561\,
            I => \row_counter.internal_count_2\
        );

    \I__667\ : InMux
    port map (
            O => \N__3558\,
            I => \row_counter.n697\
        );

    \I__666\ : InMux
    port map (
            O => \N__3555\,
            I => \N__3552\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__3552\,
            I => \N__3548\
        );

    \I__664\ : InMux
    port map (
            O => \N__3551\,
            I => \N__3545\
        );

    \I__663\ : Odrv4
    port map (
            O => \N__3548\,
            I => \row_counter.internal_count_3\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__3545\,
            I => \row_counter.internal_count_3\
        );

    \I__661\ : InMux
    port map (
            O => \N__3540\,
            I => \row_counter.n698\
        );

    \I__660\ : InMux
    port map (
            O => \N__3537\,
            I => \N__3533\
        );

    \I__659\ : InMux
    port map (
            O => \N__3536\,
            I => \N__3530\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__3533\,
            I => \row_counter.internal_count_4\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__3530\,
            I => \row_counter.internal_count_4\
        );

    \I__656\ : InMux
    port map (
            O => \N__3525\,
            I => \N__3522\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__3522\,
            I => \N__3519\
        );

    \I__654\ : Odrv4
    port map (
            O => \N__3519\,
            I => sr_row_data_4
        );

    \I__653\ : InMux
    port map (
            O => \N__3516\,
            I => \row_counter.n699\
        );

    \I__652\ : InMux
    port map (
            O => \N__3513\,
            I => \N__3509\
        );

    \I__651\ : InMux
    port map (
            O => \N__3512\,
            I => \N__3506\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__3509\,
            I => \row_counter.internal_count_5\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__3506\,
            I => \row_counter.internal_count_5\
        );

    \I__648\ : InMux
    port map (
            O => \N__3501\,
            I => \row_counter.n700\
        );

    \I__647\ : InMux
    port map (
            O => \N__3498\,
            I => \N__3494\
        );

    \I__646\ : InMux
    port map (
            O => \N__3497\,
            I => \N__3491\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__3494\,
            I => \row_counter.internal_count_6\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__3491\,
            I => \row_counter.internal_count_6\
        );

    \I__643\ : InMux
    port map (
            O => \N__3486\,
            I => \row_counter.n701\
        );

    \I__642\ : InMux
    port map (
            O => \N__3483\,
            I => \N__3479\
        );

    \I__641\ : InMux
    port map (
            O => \N__3482\,
            I => \N__3476\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__3479\,
            I => \row_counter.internal_count_7\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__3476\,
            I => \row_counter.internal_count_7\
        );

    \I__638\ : CascadeMux
    port map (
            O => \N__3471\,
            I => \N__3468\
        );

    \I__637\ : InMux
    port map (
            O => \N__3468\,
            I => \N__3465\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__3465\,
            I => \N__3462\
        );

    \I__635\ : Odrv4
    port map (
            O => \N__3462\,
            I => sr_row_data_7
        );

    \I__634\ : InMux
    port map (
            O => \N__3459\,
            I => \row_counter.n702\
        );

    \I__633\ : InMux
    port map (
            O => \N__3456\,
            I => \N__3453\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__3453\,
            I => \N__3450\
        );

    \I__631\ : Span4Mux_h
    port map (
            O => \N__3450\,
            I => \N__3447\
        );

    \I__630\ : Sp12to4
    port map (
            O => \N__3447\,
            I => \N__3444\
        );

    \I__629\ : Span12Mux_v
    port map (
            O => \N__3444\,
            I => \N__3441\
        );

    \I__628\ : Odrv12
    port map (
            O => \N__3441\,
            I => en_rowpack_c
        );

    \I__627\ : CEMux
    port map (
            O => \N__3438\,
            I => \N__3434\
        );

    \I__626\ : CEMux
    port map (
            O => \N__3437\,
            I => \N__3431\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__3434\,
            I => \N__3428\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__3431\,
            I => \N__3425\
        );

    \I__623\ : Odrv12
    port map (
            O => \N__3428\,
            I => n189
        );

    \I__622\ : Odrv4
    port map (
            O => \N__3425\,
            I => n189
        );

    \I__621\ : InMux
    port map (
            O => \N__3420\,
            I => \N__3417\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__3417\,
            I => \N__3413\
        );

    \I__619\ : InMux
    port map (
            O => \N__3416\,
            I => \N__3410\
        );

    \I__618\ : Span4Mux_v
    port map (
            O => \N__3413\,
            I => \N__3405\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__3410\,
            I => \N__3405\
        );

    \I__616\ : Span4Mux_v
    port map (
            O => \N__3405\,
            I => \N__3402\
        );

    \I__615\ : Span4Mux_v
    port map (
            O => \N__3402\,
            I => \N__3399\
        );

    \I__614\ : Sp12to4
    port map (
            O => \N__3399\,
            I => \N__3396\
        );

    \I__613\ : Odrv12
    port map (
            O => \N__3396\,
            I => sr_data_c
        );

    \I__612\ : InMux
    port map (
            O => \N__3393\,
            I => \N__3390\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__3390\,
            I => \N__3385\
        );

    \I__610\ : InMux
    port map (
            O => \N__3389\,
            I => \N__3380\
        );

    \I__609\ : InMux
    port map (
            O => \N__3388\,
            I => \N__3380\
        );

    \I__608\ : Odrv4
    port map (
            O => \N__3385\,
            I => shifted_data_0
        );

    \I__607\ : LocalMux
    port map (
            O => \N__3380\,
            I => shifted_data_0
        );

    \I__606\ : InMux
    port map (
            O => \N__3375\,
            I => \N__3371\
        );

    \I__605\ : CascadeMux
    port map (
            O => \N__3374\,
            I => \N__3368\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__3371\,
            I => \N__3364\
        );

    \I__603\ : InMux
    port map (
            O => \N__3368\,
            I => \N__3361\
        );

    \I__602\ : InMux
    port map (
            O => \N__3367\,
            I => \N__3358\
        );

    \I__601\ : Odrv4
    port map (
            O => \N__3364\,
            I => shifted_data_1
        );

    \I__600\ : LocalMux
    port map (
            O => \N__3361\,
            I => shifted_data_1
        );

    \I__599\ : LocalMux
    port map (
            O => \N__3358\,
            I => shifted_data_1
        );

    \I__598\ : CascadeMux
    port map (
            O => \N__3351\,
            I => \N__3347\
        );

    \I__597\ : InMux
    port map (
            O => \N__3350\,
            I => \N__3344\
        );

    \I__596\ : InMux
    port map (
            O => \N__3347\,
            I => \N__3340\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__3344\,
            I => \N__3337\
        );

    \I__594\ : InMux
    port map (
            O => \N__3343\,
            I => \N__3334\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__3340\,
            I => \N__3331\
        );

    \I__592\ : Odrv12
    port map (
            O => \N__3337\,
            I => shifted_data_2
        );

    \I__591\ : LocalMux
    port map (
            O => \N__3334\,
            I => shifted_data_2
        );

    \I__590\ : Odrv4
    port map (
            O => \N__3331\,
            I => shifted_data_2
        );

    \I__589\ : InMux
    port map (
            O => \N__3324\,
            I => \N__3321\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__3321\,
            I => \N__3312\
        );

    \I__587\ : InMux
    port map (
            O => \N__3320\,
            I => \N__3303\
        );

    \I__586\ : InMux
    port map (
            O => \N__3319\,
            I => \N__3303\
        );

    \I__585\ : InMux
    port map (
            O => \N__3318\,
            I => \N__3303\
        );

    \I__584\ : InMux
    port map (
            O => \N__3317\,
            I => \N__3303\
        );

    \I__583\ : CascadeMux
    port map (
            O => \N__3316\,
            I => \N__3299\
        );

    \I__582\ : CascadeMux
    port map (
            O => \N__3315\,
            I => \N__3291\
        );

    \I__581\ : Span4Mux_v
    port map (
            O => \N__3312\,
            I => \N__3286\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__3303\,
            I => \N__3283\
        );

    \I__579\ : InMux
    port map (
            O => \N__3302\,
            I => \N__3270\
        );

    \I__578\ : InMux
    port map (
            O => \N__3299\,
            I => \N__3270\
        );

    \I__577\ : InMux
    port map (
            O => \N__3298\,
            I => \N__3270\
        );

    \I__576\ : InMux
    port map (
            O => \N__3297\,
            I => \N__3270\
        );

    \I__575\ : InMux
    port map (
            O => \N__3296\,
            I => \N__3270\
        );

    \I__574\ : InMux
    port map (
            O => \N__3295\,
            I => \N__3270\
        );

    \I__573\ : InMux
    port map (
            O => \N__3294\,
            I => \N__3261\
        );

    \I__572\ : InMux
    port map (
            O => \N__3291\,
            I => \N__3261\
        );

    \I__571\ : InMux
    port map (
            O => \N__3290\,
            I => \N__3261\
        );

    \I__570\ : InMux
    port map (
            O => \N__3289\,
            I => \N__3261\
        );

    \I__569\ : Odrv4
    port map (
            O => \N__3286\,
            I => n330
        );

    \I__568\ : Odrv12
    port map (
            O => \N__3283\,
            I => n330
        );

    \I__567\ : LocalMux
    port map (
            O => \N__3270\,
            I => n330
        );

    \I__566\ : LocalMux
    port map (
            O => \N__3261\,
            I => n330
        );

    \I__565\ : CascadeMux
    port map (
            O => \N__3252\,
            I => \N__3249\
        );

    \I__564\ : InMux
    port map (
            O => \N__3249\,
            I => \N__3245\
        );

    \I__563\ : CascadeMux
    port map (
            O => \N__3248\,
            I => \N__3239\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__3245\,
            I => \N__3233\
        );

    \I__561\ : InMux
    port map (
            O => \N__3244\,
            I => \N__3228\
        );

    \I__560\ : InMux
    port map (
            O => \N__3243\,
            I => \N__3228\
        );

    \I__559\ : InMux
    port map (
            O => \N__3242\,
            I => \N__3223\
        );

    \I__558\ : InMux
    port map (
            O => \N__3239\,
            I => \N__3223\
        );

    \I__557\ : CascadeMux
    port map (
            O => \N__3238\,
            I => \N__3217\
        );

    \I__556\ : CascadeMux
    port map (
            O => \N__3237\,
            I => \N__3213\
        );

    \I__555\ : CascadeMux
    port map (
            O => \N__3236\,
            I => \N__3207\
        );

    \I__554\ : Span4Mux_v
    port map (
            O => \N__3233\,
            I => \N__3204\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__3228\,
            I => \N__3199\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__3223\,
            I => \N__3199\
        );

    \I__551\ : InMux
    port map (
            O => \N__3222\,
            I => \N__3186\
        );

    \I__550\ : InMux
    port map (
            O => \N__3221\,
            I => \N__3186\
        );

    \I__549\ : InMux
    port map (
            O => \N__3220\,
            I => \N__3186\
        );

    \I__548\ : InMux
    port map (
            O => \N__3217\,
            I => \N__3186\
        );

    \I__547\ : InMux
    port map (
            O => \N__3216\,
            I => \N__3186\
        );

    \I__546\ : InMux
    port map (
            O => \N__3213\,
            I => \N__3186\
        );

    \I__545\ : InMux
    port map (
            O => \N__3212\,
            I => \N__3183\
        );

    \I__544\ : InMux
    port map (
            O => \N__3211\,
            I => \N__3176\
        );

    \I__543\ : InMux
    port map (
            O => \N__3210\,
            I => \N__3176\
        );

    \I__542\ : InMux
    port map (
            O => \N__3207\,
            I => \N__3176\
        );

    \I__541\ : Odrv4
    port map (
            O => \N__3204\,
            I => n169
        );

    \I__540\ : Odrv12
    port map (
            O => \N__3199\,
            I => n169
        );

    \I__539\ : LocalMux
    port map (
            O => \N__3186\,
            I => n169
        );

    \I__538\ : LocalMux
    port map (
            O => \N__3183\,
            I => n169
        );

    \I__537\ : LocalMux
    port map (
            O => \N__3176\,
            I => n169
        );

    \I__536\ : InMux
    port map (
            O => \N__3165\,
            I => \N__3161\
        );

    \I__535\ : CascadeMux
    port map (
            O => \N__3164\,
            I => \N__3157\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__3161\,
            I => \N__3154\
        );

    \I__533\ : InMux
    port map (
            O => \N__3160\,
            I => \N__3151\
        );

    \I__532\ : InMux
    port map (
            O => \N__3157\,
            I => \N__3148\
        );

    \I__531\ : Odrv4
    port map (
            O => \N__3154\,
            I => shifted_data_3
        );

    \I__530\ : LocalMux
    port map (
            O => \N__3151\,
            I => shifted_data_3
        );

    \I__529\ : LocalMux
    port map (
            O => \N__3148\,
            I => shifted_data_3
        );

    \I__528\ : CascadeMux
    port map (
            O => \N__3141\,
            I => \N__3137\
        );

    \I__527\ : InMux
    port map (
            O => \N__3140\,
            I => \N__3134\
        );

    \I__526\ : InMux
    port map (
            O => \N__3137\,
            I => \N__3130\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__3134\,
            I => \N__3127\
        );

    \I__524\ : InMux
    port map (
            O => \N__3133\,
            I => \N__3124\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__3130\,
            I => \N__3121\
        );

    \I__522\ : Odrv12
    port map (
            O => \N__3127\,
            I => shifted_data_4
        );

    \I__521\ : LocalMux
    port map (
            O => \N__3124\,
            I => shifted_data_4
        );

    \I__520\ : Odrv4
    port map (
            O => \N__3121\,
            I => shifted_data_4
        );

    \I__519\ : InMux
    port map (
            O => \N__3114\,
            I => \N__3111\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__3111\,
            I => \N__3106\
        );

    \I__517\ : InMux
    port map (
            O => \N__3110\,
            I => \N__3103\
        );

    \I__516\ : InMux
    port map (
            O => \N__3109\,
            I => \N__3100\
        );

    \I__515\ : Odrv4
    port map (
            O => \N__3106\,
            I => shifted_data_0_adj_115
        );

    \I__514\ : LocalMux
    port map (
            O => \N__3103\,
            I => shifted_data_0_adj_115
        );

    \I__513\ : LocalMux
    port map (
            O => \N__3100\,
            I => shifted_data_0_adj_115
        );

    \I__512\ : InMux
    port map (
            O => \N__3093\,
            I => \row_counter.n752\
        );

    \I__511\ : InMux
    port map (
            O => \N__3090\,
            I => \row_counter.n753\
        );

    \I__510\ : InMux
    port map (
            O => \N__3087\,
            I => \row_counter.n754\
        );

    \I__509\ : InMux
    port map (
            O => \N__3084\,
            I => \row_counter.n755\
        );

    \I__508\ : InMux
    port map (
            O => \N__3081\,
            I => \row_counter.n756\
        );

    \I__507\ : InMux
    port map (
            O => \N__3078\,
            I => \row_counter.n757\
        );

    \I__506\ : InMux
    port map (
            O => \N__3075\,
            I => \row_counter.n743\
        );

    \I__505\ : InMux
    port map (
            O => \N__3072\,
            I => \row_counter.n744\
        );

    \I__504\ : InMux
    port map (
            O => \N__3069\,
            I => \row_counter.n745\
        );

    \I__503\ : InMux
    port map (
            O => \N__3066\,
            I => \row_counter.n746\
        );

    \I__502\ : InMux
    port map (
            O => \N__3063\,
            I => \row_counter.n747\
        );

    \I__501\ : InMux
    port map (
            O => \N__3060\,
            I => \row_counter.n748\
        );

    \I__500\ : InMux
    port map (
            O => \N__3057\,
            I => \row_counter.n749\
        );

    \I__499\ : InMux
    port map (
            O => \N__3054\,
            I => \bfn_5_8_0_\
        );

    \I__498\ : InMux
    port map (
            O => \N__3051\,
            I => \row_counter.n751\
        );

    \I__497\ : CascadeMux
    port map (
            O => \N__3048\,
            I => \N__3044\
        );

    \I__496\ : InMux
    port map (
            O => \N__3047\,
            I => \N__3040\
        );

    \I__495\ : InMux
    port map (
            O => \N__3044\,
            I => \N__3037\
        );

    \I__494\ : InMux
    port map (
            O => \N__3043\,
            I => \N__3034\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__3040\,
            I => shifted_data_12
        );

    \I__492\ : LocalMux
    port map (
            O => \N__3037\,
            I => shifted_data_12
        );

    \I__491\ : LocalMux
    port map (
            O => \N__3034\,
            I => shifted_data_12
        );

    \I__490\ : InMux
    port map (
            O => \N__3027\,
            I => \N__3022\
        );

    \I__489\ : InMux
    port map (
            O => \N__3026\,
            I => \N__3017\
        );

    \I__488\ : InMux
    port map (
            O => \N__3025\,
            I => \N__3017\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__3022\,
            I => shifted_data_13
        );

    \I__486\ : LocalMux
    port map (
            O => \N__3017\,
            I => shifted_data_13
        );

    \I__485\ : InMux
    port map (
            O => \N__3012\,
            I => \N__3007\
        );

    \I__484\ : InMux
    port map (
            O => \N__3011\,
            I => \N__3002\
        );

    \I__483\ : InMux
    port map (
            O => \N__3010\,
            I => \N__3002\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__3007\,
            I => shifted_data_8
        );

    \I__481\ : LocalMux
    port map (
            O => \N__3002\,
            I => shifted_data_8
        );

    \I__480\ : CascadeMux
    port map (
            O => \N__2997\,
            I => \N__2993\
        );

    \I__479\ : InMux
    port map (
            O => \N__2996\,
            I => \N__2989\
        );

    \I__478\ : InMux
    port map (
            O => \N__2993\,
            I => \N__2986\
        );

    \I__477\ : InMux
    port map (
            O => \N__2992\,
            I => \N__2983\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__2989\,
            I => shifted_data_9
        );

    \I__475\ : LocalMux
    port map (
            O => \N__2986\,
            I => shifted_data_9
        );

    \I__474\ : LocalMux
    port map (
            O => \N__2983\,
            I => shifted_data_9
        );

    \I__473\ : InMux
    port map (
            O => \N__2976\,
            I => \N__2971\
        );

    \I__472\ : InMux
    port map (
            O => \N__2975\,
            I => \N__2968\
        );

    \I__471\ : InMux
    port map (
            O => \N__2974\,
            I => \N__2965\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__2971\,
            I => shifted_data_10
        );

    \I__469\ : LocalMux
    port map (
            O => \N__2968\,
            I => shifted_data_10
        );

    \I__468\ : LocalMux
    port map (
            O => \N__2965\,
            I => shifted_data_10
        );

    \I__467\ : InMux
    port map (
            O => \N__2958\,
            I => \N__2953\
        );

    \I__466\ : InMux
    port map (
            O => \N__2957\,
            I => \N__2948\
        );

    \I__465\ : InMux
    port map (
            O => \N__2956\,
            I => \N__2948\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__2953\,
            I => shifted_data_5
        );

    \I__463\ : LocalMux
    port map (
            O => \N__2948\,
            I => shifted_data_5
        );

    \I__462\ : InMux
    port map (
            O => \N__2943\,
            I => \N__2938\
        );

    \I__461\ : InMux
    port map (
            O => \N__2942\,
            I => \N__2933\
        );

    \I__460\ : InMux
    port map (
            O => \N__2941\,
            I => \N__2933\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__2938\,
            I => shifted_data_6
        );

    \I__458\ : LocalMux
    port map (
            O => \N__2933\,
            I => shifted_data_6
        );

    \I__457\ : CascadeMux
    port map (
            O => \N__2928\,
            I => \N__2924\
        );

    \I__456\ : InMux
    port map (
            O => \N__2927\,
            I => \N__2920\
        );

    \I__455\ : InMux
    port map (
            O => \N__2924\,
            I => \N__2917\
        );

    \I__454\ : InMux
    port map (
            O => \N__2923\,
            I => \N__2914\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__2920\,
            I => shifted_data_7
        );

    \I__452\ : LocalMux
    port map (
            O => \N__2917\,
            I => shifted_data_7
        );

    \I__451\ : LocalMux
    port map (
            O => \N__2914\,
            I => shifted_data_7
        );

    \I__450\ : InMux
    port map (
            O => \N__2907\,
            I => \bfn_5_7_0_\
        );

    \I__449\ : InMux
    port map (
            O => \N__2904\,
            I => \N__2901\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__2901\,
            I => n2_adj_99
        );

    \I__447\ : InMux
    port map (
            O => \N__2898\,
            I => \N__2895\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__2895\,
            I => n11
        );

    \I__445\ : CascadeMux
    port map (
            O => \N__2892\,
            I => \n823_cascade_\
        );

    \I__444\ : InMux
    port map (
            O => \N__2889\,
            I => \N__2886\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__2886\,
            I => n781
        );

    \I__442\ : InMux
    port map (
            O => \N__2883\,
            I => \N__2880\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__2880\,
            I => n827
        );

    \I__440\ : InMux
    port map (
            O => \N__2877\,
            I => \N__2871\
        );

    \I__439\ : InMux
    port map (
            O => \N__2876\,
            I => \N__2871\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__2871\,
            I => \N__2868\
        );

    \I__437\ : Span4Mux_v
    port map (
            O => \N__2868\,
            I => \N__2865\
        );

    \I__436\ : Sp12to4
    port map (
            O => \N__2865\,
            I => \N__2862\
        );

    \I__435\ : Odrv12
    port map (
            O => \N__2862\,
            I => sr_sel_row_c
        );

    \I__434\ : CascadeMux
    port map (
            O => \N__2859\,
            I => \n169_cascade_\
        );

    \I__433\ : InMux
    port map (
            O => \N__2856\,
            I => \N__2850\
        );

    \I__432\ : InMux
    port map (
            O => \N__2855\,
            I => \N__2850\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__2850\,
            I => \N__2847\
        );

    \I__430\ : Span12Mux_h
    port map (
            O => \N__2847\,
            I => \N__2844\
        );

    \I__429\ : Span12Mux_v
    port map (
            O => \N__2844\,
            I => \N__2841\
        );

    \I__428\ : Odrv12
    port map (
            O => \N__2841\,
            I => sr_sel_div_c
        );

    \I__427\ : InMux
    port map (
            O => \N__2838\,
            I => \N__2830\
        );

    \I__426\ : InMux
    port map (
            O => \N__2837\,
            I => \N__2830\
        );

    \I__425\ : InMux
    port map (
            O => \N__2836\,
            I => \N__2825\
        );

    \I__424\ : InMux
    port map (
            O => \N__2835\,
            I => \N__2825\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__2830\,
            I => \N__2820\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__2825\,
            I => \N__2820\
        );

    \I__421\ : Span4Mux_v
    port map (
            O => \N__2820\,
            I => \N__2817\
        );

    \I__420\ : Sp12to4
    port map (
            O => \N__2817\,
            I => \N__2814\
        );

    \I__419\ : Odrv12
    port map (
            O => \N__2814\,
            I => sr_reset_c
        );

    \I__418\ : CascadeMux
    port map (
            O => \N__2811\,
            I => \n330_cascade_\
        );

    \I__417\ : InMux
    port map (
            O => \N__2808\,
            I => \N__2803\
        );

    \I__416\ : InMux
    port map (
            O => \N__2807\,
            I => \N__2798\
        );

    \I__415\ : InMux
    port map (
            O => \N__2806\,
            I => \N__2798\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__2803\,
            I => shifted_data_14
        );

    \I__413\ : LocalMux
    port map (
            O => \N__2798\,
            I => shifted_data_14
        );

    \I__412\ : InMux
    port map (
            O => \N__2793\,
            I => \N__2789\
        );

    \I__411\ : InMux
    port map (
            O => \N__2792\,
            I => \N__2786\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__2789\,
            I => shifted_data_15
        );

    \I__409\ : LocalMux
    port map (
            O => \N__2786\,
            I => shifted_data_15
        );

    \I__408\ : InMux
    port map (
            O => \N__2781\,
            I => \N__2776\
        );

    \I__407\ : InMux
    port map (
            O => \N__2780\,
            I => \N__2771\
        );

    \I__406\ : InMux
    port map (
            O => \N__2779\,
            I => \N__2771\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__2776\,
            I => shifted_data_11
        );

    \I__404\ : LocalMux
    port map (
            O => \N__2771\,
            I => shifted_data_11
        );

    \I__403\ : InMux
    port map (
            O => \N__2766\,
            I => \N__2763\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__2763\,
            I => \N__2760\
        );

    \I__401\ : Odrv4
    port map (
            O => \N__2760\,
            I => sr_divider_data_10
        );

    \I__400\ : InMux
    port map (
            O => \N__2757\,
            I => \N__2754\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__2754\,
            I => \N__2751\
        );

    \I__398\ : Odrv12
    port map (
            O => \N__2751\,
            I => sr_divider_data_6
        );

    \I__397\ : InMux
    port map (
            O => \N__2748\,
            I => \N__2745\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__2745\,
            I => \N__2742\
        );

    \I__395\ : Odrv4
    port map (
            O => \N__2742\,
            I => sr_divider_data_9
        );

    \I__394\ : CascadeMux
    port map (
            O => \N__2739\,
            I => \N__2736\
        );

    \I__393\ : InMux
    port map (
            O => \N__2736\,
            I => \N__2733\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__2733\,
            I => \N__2730\
        );

    \I__391\ : Odrv12
    port map (
            O => \N__2730\,
            I => sr_divider_data_4
        );

    \I__390\ : InMux
    port map (
            O => \N__2727\,
            I => \N__2724\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__2724\,
            I => \N__2721\
        );

    \I__388\ : Odrv12
    port map (
            O => \N__2721\,
            I => sr_divider_data_5
        );

    \I__387\ : InMux
    port map (
            O => \N__2718\,
            I => \N__2715\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__2715\,
            I => \N__2712\
        );

    \I__385\ : Span4Mux_v
    port map (
            O => \N__2712\,
            I => \N__2709\
        );

    \I__384\ : Odrv4
    port map (
            O => \N__2709\,
            I => sr_divider_data_8
        );

    \I__383\ : InMux
    port map (
            O => \N__2706\,
            I => \N__2703\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__2703\,
            I => \N__2700\
        );

    \I__381\ : Odrv12
    port map (
            O => \N__2700\,
            I => sr_divider_data_7
        );

    \I__380\ : InMux
    port map (
            O => \N__2697\,
            I => \N__2694\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__2694\,
            I => n8
        );

    \I__378\ : InMux
    port map (
            O => \N__2691\,
            I => \N__2688\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__2688\,
            I => n3_adj_118
        );

    \I__376\ : InMux
    port map (
            O => \N__2685\,
            I => \N__2682\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__2682\,
            I => n15
        );

    \I__374\ : InMux
    port map (
            O => \N__2679\,
            I => \N__2676\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__2676\,
            I => n7
        );

    \I__372\ : CascadeMux
    port map (
            O => \N__2673\,
            I => \N__2670\
        );

    \I__371\ : InMux
    port map (
            O => \N__2670\,
            I => \N__2667\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__2667\,
            I => n10
        );

    \I__369\ : InMux
    port map (
            O => \N__2664\,
            I => \N__2661\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__2661\,
            I => n14
        );

    \I__367\ : CascadeMux
    port map (
            O => \N__2658\,
            I => \N__2655\
        );

    \I__366\ : InMux
    port map (
            O => \N__2655\,
            I => \N__2652\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__2652\,
            I => sr_divider_data_13
        );

    \I__364\ : InMux
    port map (
            O => \N__2649\,
            I => \N__2641\
        );

    \I__363\ : InMux
    port map (
            O => \N__2648\,
            I => \N__2641\
        );

    \I__362\ : InMux
    port map (
            O => \N__2647\,
            I => \N__2636\
        );

    \I__361\ : InMux
    port map (
            O => \N__2646\,
            I => \N__2636\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__2641\,
            I => count_done
        );

    \I__359\ : LocalMux
    port map (
            O => \N__2636\,
            I => count_done
        );

    \I__358\ : ClkMux
    port map (
            O => \N__2631\,
            I => \N__2619\
        );

    \I__357\ : ClkMux
    port map (
            O => \N__2630\,
            I => \N__2619\
        );

    \I__356\ : ClkMux
    port map (
            O => \N__2629\,
            I => \N__2619\
        );

    \I__355\ : ClkMux
    port map (
            O => \N__2628\,
            I => \N__2619\
        );

    \I__354\ : GlobalMux
    port map (
            O => \N__2619\,
            I => \N__2616\
        );

    \I__353\ : gio2CtrlBuf
    port map (
            O => \N__2616\,
            I => laser_pulse_c
        );

    \I__352\ : CascadeMux
    port map (
            O => \N__2613\,
            I => \N__2610\
        );

    \I__351\ : InMux
    port map (
            O => \N__2610\,
            I => \N__2607\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__2607\,
            I => \N__2604\
        );

    \I__349\ : Odrv12
    port map (
            O => \N__2604\,
            I => sr_divider_data_2
        );

    \I__348\ : CascadeMux
    port map (
            O => \N__2601\,
            I => \N__2598\
        );

    \I__347\ : InMux
    port map (
            O => \N__2598\,
            I => \N__2595\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__2595\,
            I => \N__2592\
        );

    \I__345\ : Odrv12
    port map (
            O => \N__2592\,
            I => sr_divider_data_14
        );

    \I__344\ : CascadeMux
    port map (
            O => \N__2589\,
            I => \N__2586\
        );

    \I__343\ : InMux
    port map (
            O => \N__2586\,
            I => \N__2583\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__2583\,
            I => \N__2580\
        );

    \I__341\ : Odrv4
    port map (
            O => \N__2580\,
            I => sr_divider_data_15
        );

    \I__340\ : InMux
    port map (
            O => \N__2577\,
            I => \N__2574\
        );

    \I__339\ : LocalMux
    port map (
            O => \N__2574\,
            I => \N__2571\
        );

    \I__338\ : Odrv4
    port map (
            O => \N__2571\,
            I => sr_divider_data_0
        );

    \I__337\ : InMux
    port map (
            O => \N__2568\,
            I => \N__2565\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__2565\,
            I => \N__2562\
        );

    \I__335\ : Odrv4
    port map (
            O => \N__2562\,
            I => sr_divider_data_3
        );

    \I__334\ : InMux
    port map (
            O => \N__2559\,
            I => \N__2556\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__2556\,
            I => \N__2553\
        );

    \I__332\ : Odrv4
    port map (
            O => \N__2553\,
            I => sr_divider_data_12
        );

    \I__331\ : InMux
    port map (
            O => \N__2550\,
            I => \N__2547\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__2547\,
            I => \N__2544\
        );

    \I__329\ : Odrv12
    port map (
            O => \N__2544\,
            I => sr_divider_data_1
        );

    \I__328\ : InMux
    port map (
            O => \N__2541\,
            I => \N__2537\
        );

    \I__327\ : InMux
    port map (
            O => \N__2540\,
            I => \N__2534\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__2537\,
            I => \N__2531\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__2534\,
            I => \pulse_counter.internal_count_14\
        );

    \I__324\ : Odrv4
    port map (
            O => \N__2531\,
            I => \pulse_counter.internal_count_14\
        );

    \I__323\ : InMux
    port map (
            O => \N__2526\,
            I => \pulse_counter.n725\
        );

    \I__322\ : InMux
    port map (
            O => \N__2523\,
            I => \N__2519\
        );

    \I__321\ : InMux
    port map (
            O => \N__2522\,
            I => \N__2516\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__2519\,
            I => \N__2513\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__2516\,
            I => \pulse_counter.internal_count_15\
        );

    \I__318\ : Odrv4
    port map (
            O => \N__2513\,
            I => \pulse_counter.internal_count_15\
        );

    \I__317\ : InMux
    port map (
            O => \N__2508\,
            I => \pulse_counter.n726\
        );

    \I__316\ : InMux
    port map (
            O => \N__2505\,
            I => \N__2502\
        );

    \I__315\ : LocalMux
    port map (
            O => \N__2502\,
            I => \pulse_counter.n13\
        );

    \I__314\ : InMux
    port map (
            O => \N__2499\,
            I => \bfn_2_9_0_\
        );

    \I__313\ : InMux
    port map (
            O => \N__2496\,
            I => \N__2493\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__2493\,
            I => \N__2490\
        );

    \I__311\ : Odrv4
    port map (
            O => \N__2490\,
            I => n4_adj_116
        );

    \I__310\ : InMux
    port map (
            O => \N__2487\,
            I => \N__2484\
        );

    \I__309\ : LocalMux
    port map (
            O => \N__2484\,
            I => \N__2481\
        );

    \I__308\ : Odrv4
    port map (
            O => \N__2481\,
            I => n5_adj_120
        );

    \I__307\ : InMux
    port map (
            O => \N__2478\,
            I => \N__2475\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__2475\,
            I => \N__2472\
        );

    \I__305\ : Odrv4
    port map (
            O => \N__2472\,
            I => n1_adj_117
        );

    \I__304\ : InMux
    port map (
            O => \N__2469\,
            I => \N__2466\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__2466\,
            I => n9
        );

    \I__302\ : CascadeMux
    port map (
            O => \N__2463\,
            I => \n795_cascade_\
        );

    \I__301\ : InMux
    port map (
            O => \N__2460\,
            I => \N__2457\
        );

    \I__300\ : LocalMux
    port map (
            O => \N__2457\,
            I => \N__2454\
        );

    \I__299\ : Odrv4
    port map (
            O => \N__2454\,
            I => n6_adj_119
        );

    \I__298\ : InMux
    port map (
            O => \N__2451\,
            I => \N__2448\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__2448\,
            I => n12
        );

    \I__296\ : InMux
    port map (
            O => \N__2445\,
            I => \N__2442\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__2442\,
            I => n16
        );

    \I__294\ : CascadeMux
    port map (
            O => \N__2439\,
            I => \n817_cascade_\
        );

    \I__293\ : InMux
    port map (
            O => \N__2436\,
            I => \N__2433\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__2433\,
            I => n787
        );

    \I__291\ : CascadeMux
    port map (
            O => \N__2430\,
            I => \n825_cascade_\
        );

    \I__290\ : InMux
    port map (
            O => \N__2427\,
            I => \N__2424\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__2424\,
            I => sr_divider_data_11
        );

    \I__288\ : InMux
    port map (
            O => \N__2421\,
            I => \N__2417\
        );

    \I__287\ : InMux
    port map (
            O => \N__2420\,
            I => \N__2414\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__2417\,
            I => \pulse_counter.internal_count_5\
        );

    \I__285\ : LocalMux
    port map (
            O => \N__2414\,
            I => \pulse_counter.internal_count_5\
        );

    \I__284\ : InMux
    port map (
            O => \N__2409\,
            I => \pulse_counter.n716\
        );

    \I__283\ : InMux
    port map (
            O => \N__2406\,
            I => \N__2402\
        );

    \I__282\ : InMux
    port map (
            O => \N__2405\,
            I => \N__2399\
        );

    \I__281\ : LocalMux
    port map (
            O => \N__2402\,
            I => \pulse_counter.internal_count_6\
        );

    \I__280\ : LocalMux
    port map (
            O => \N__2399\,
            I => \pulse_counter.internal_count_6\
        );

    \I__279\ : InMux
    port map (
            O => \N__2394\,
            I => \pulse_counter.n717\
        );

    \I__278\ : InMux
    port map (
            O => \N__2391\,
            I => \N__2387\
        );

    \I__277\ : InMux
    port map (
            O => \N__2390\,
            I => \N__2384\
        );

    \I__276\ : LocalMux
    port map (
            O => \N__2387\,
            I => \pulse_counter.internal_count_7\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__2384\,
            I => \pulse_counter.internal_count_7\
        );

    \I__274\ : InMux
    port map (
            O => \N__2379\,
            I => \pulse_counter.n718\
        );

    \I__273\ : InMux
    port map (
            O => \N__2376\,
            I => \N__2372\
        );

    \I__272\ : InMux
    port map (
            O => \N__2375\,
            I => \N__2369\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__2372\,
            I => \pulse_counter.internal_count_8\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__2369\,
            I => \pulse_counter.internal_count_8\
        );

    \I__269\ : InMux
    port map (
            O => \N__2364\,
            I => \bfn_2_8_0_\
        );

    \I__268\ : InMux
    port map (
            O => \N__2361\,
            I => \N__2357\
        );

    \I__267\ : InMux
    port map (
            O => \N__2360\,
            I => \N__2354\
        );

    \I__266\ : LocalMux
    port map (
            O => \N__2357\,
            I => \pulse_counter.internal_count_9\
        );

    \I__265\ : LocalMux
    port map (
            O => \N__2354\,
            I => \pulse_counter.internal_count_9\
        );

    \I__264\ : InMux
    port map (
            O => \N__2349\,
            I => \pulse_counter.n720\
        );

    \I__263\ : InMux
    port map (
            O => \N__2346\,
            I => \N__2342\
        );

    \I__262\ : InMux
    port map (
            O => \N__2345\,
            I => \N__2339\
        );

    \I__261\ : LocalMux
    port map (
            O => \N__2342\,
            I => \pulse_counter.internal_count_10\
        );

    \I__260\ : LocalMux
    port map (
            O => \N__2339\,
            I => \pulse_counter.internal_count_10\
        );

    \I__259\ : InMux
    port map (
            O => \N__2334\,
            I => \pulse_counter.n721\
        );

    \I__258\ : InMux
    port map (
            O => \N__2331\,
            I => \N__2327\
        );

    \I__257\ : InMux
    port map (
            O => \N__2330\,
            I => \N__2324\
        );

    \I__256\ : LocalMux
    port map (
            O => \N__2327\,
            I => \pulse_counter.internal_count_11\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__2324\,
            I => \pulse_counter.internal_count_11\
        );

    \I__254\ : InMux
    port map (
            O => \N__2319\,
            I => \pulse_counter.n722\
        );

    \I__253\ : InMux
    port map (
            O => \N__2316\,
            I => \N__2312\
        );

    \I__252\ : InMux
    port map (
            O => \N__2315\,
            I => \N__2309\
        );

    \I__251\ : LocalMux
    port map (
            O => \N__2312\,
            I => \pulse_counter.internal_count_12\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__2309\,
            I => \pulse_counter.internal_count_12\
        );

    \I__249\ : InMux
    port map (
            O => \N__2304\,
            I => \pulse_counter.n723\
        );

    \I__248\ : InMux
    port map (
            O => \N__2301\,
            I => \N__2297\
        );

    \I__247\ : InMux
    port map (
            O => \N__2300\,
            I => \N__2294\
        );

    \I__246\ : LocalMux
    port map (
            O => \N__2297\,
            I => \pulse_counter.internal_count_13\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__2294\,
            I => \pulse_counter.internal_count_13\
        );

    \I__244\ : InMux
    port map (
            O => \N__2289\,
            I => \pulse_counter.n724\
        );

    \I__243\ : CascadeMux
    port map (
            O => \N__2286\,
            I => \N__2283\
        );

    \I__242\ : InMux
    port map (
            O => \N__2283\,
            I => \N__2277\
        );

    \I__241\ : InMux
    port map (
            O => \N__2282\,
            I => \N__2277\
        );

    \I__240\ : LocalMux
    port map (
            O => \N__2277\,
            I => \N__2274\
        );

    \I__239\ : Span12Mux_h
    port map (
            O => \N__2274\,
            I => \N__2271\
        );

    \I__238\ : Span12Mux_v
    port map (
            O => \N__2271\,
            I => \N__2268\
        );

    \I__237\ : Odrv12
    port map (
            O => \N__2268\,
            I => divide_enable_c
        );

    \I__236\ : CEMux
    port map (
            O => \N__2265\,
            I => \N__2262\
        );

    \I__235\ : LocalMux
    port map (
            O => \N__2262\,
            I => \N__2258\
        );

    \I__234\ : CEMux
    port map (
            O => \N__2261\,
            I => \N__2255\
        );

    \I__233\ : Span4Mux_v
    port map (
            O => \N__2258\,
            I => \N__2250\
        );

    \I__232\ : LocalMux
    port map (
            O => \N__2255\,
            I => \N__2250\
        );

    \I__231\ : Span4Mux_h
    port map (
            O => \N__2250\,
            I => \N__2247\
        );

    \I__230\ : Odrv4
    port map (
            O => \N__2247\,
            I => n176
        );

    \I__229\ : InMux
    port map (
            O => \N__2244\,
            I => \N__2240\
        );

    \I__228\ : InMux
    port map (
            O => \N__2243\,
            I => \N__2237\
        );

    \I__227\ : LocalMux
    port map (
            O => \N__2240\,
            I => output_state
        );

    \I__226\ : LocalMux
    port map (
            O => \N__2237\,
            I => output_state
        );

    \I__225\ : InMux
    port map (
            O => \N__2232\,
            I => \N__2229\
        );

    \I__224\ : LocalMux
    port map (
            O => \N__2229\,
            I => \N__2226\
        );

    \I__223\ : Span4Mux_v
    port map (
            O => \N__2226\,
            I => \N__2223\
        );

    \I__222\ : Span4Mux_v
    port map (
            O => \N__2223\,
            I => \N__2220\
        );

    \I__221\ : Sp12to4
    port map (
            O => \N__2220\,
            I => \N__2217\
        );

    \I__220\ : Odrv12
    port map (
            O => \N__2217\,
            I => constant_v_c
        );

    \I__219\ : InMux
    port map (
            O => \N__2214\,
            I => \N__2210\
        );

    \I__218\ : InMux
    port map (
            O => \N__2213\,
            I => \N__2207\
        );

    \I__217\ : LocalMux
    port map (
            O => \N__2210\,
            I => \pulse_counter.internal_count_0\
        );

    \I__216\ : LocalMux
    port map (
            O => \N__2207\,
            I => \pulse_counter.internal_count_0\
        );

    \I__215\ : InMux
    port map (
            O => \N__2202\,
            I => \bfn_2_7_0_\
        );

    \I__214\ : InMux
    port map (
            O => \N__2199\,
            I => \N__2195\
        );

    \I__213\ : InMux
    port map (
            O => \N__2198\,
            I => \N__2192\
        );

    \I__212\ : LocalMux
    port map (
            O => \N__2195\,
            I => \pulse_counter.internal_count_1\
        );

    \I__211\ : LocalMux
    port map (
            O => \N__2192\,
            I => \pulse_counter.internal_count_1\
        );

    \I__210\ : InMux
    port map (
            O => \N__2187\,
            I => \pulse_counter.n712\
        );

    \I__209\ : InMux
    port map (
            O => \N__2184\,
            I => \N__2180\
        );

    \I__208\ : InMux
    port map (
            O => \N__2183\,
            I => \N__2177\
        );

    \I__207\ : LocalMux
    port map (
            O => \N__2180\,
            I => \pulse_counter.internal_count_2\
        );

    \I__206\ : LocalMux
    port map (
            O => \N__2177\,
            I => \pulse_counter.internal_count_2\
        );

    \I__205\ : InMux
    port map (
            O => \N__2172\,
            I => \pulse_counter.n713\
        );

    \I__204\ : InMux
    port map (
            O => \N__2169\,
            I => \N__2165\
        );

    \I__203\ : InMux
    port map (
            O => \N__2168\,
            I => \N__2162\
        );

    \I__202\ : LocalMux
    port map (
            O => \N__2165\,
            I => \pulse_counter.internal_count_3\
        );

    \I__201\ : LocalMux
    port map (
            O => \N__2162\,
            I => \pulse_counter.internal_count_3\
        );

    \I__200\ : InMux
    port map (
            O => \N__2157\,
            I => \pulse_counter.n714\
        );

    \I__199\ : InMux
    port map (
            O => \N__2154\,
            I => \N__2150\
        );

    \I__198\ : InMux
    port map (
            O => \N__2153\,
            I => \N__2147\
        );

    \I__197\ : LocalMux
    port map (
            O => \N__2150\,
            I => \pulse_counter.internal_count_4\
        );

    \I__196\ : LocalMux
    port map (
            O => \N__2147\,
            I => \pulse_counter.internal_count_4\
        );

    \I__195\ : InMux
    port map (
            O => \N__2142\,
            I => \pulse_counter.n715\
        );

    \I__194\ : InMux
    port map (
            O => \N__2139\,
            I => \pulse_counter.n734\
        );

    \I__193\ : InMux
    port map (
            O => \N__2136\,
            I => \bfn_1_8_0_\
        );

    \I__192\ : InMux
    port map (
            O => \N__2133\,
            I => \pulse_counter.n736\
        );

    \I__191\ : InMux
    port map (
            O => \N__2130\,
            I => \pulse_counter.n737\
        );

    \I__190\ : InMux
    port map (
            O => \N__2127\,
            I => \pulse_counter.n738\
        );

    \I__189\ : InMux
    port map (
            O => \N__2124\,
            I => \pulse_counter.n739\
        );

    \I__188\ : InMux
    port map (
            O => \N__2121\,
            I => \pulse_counter.n740\
        );

    \I__187\ : InMux
    port map (
            O => \N__2118\,
            I => \pulse_counter.n741\
        );

    \I__186\ : InMux
    port map (
            O => \N__2115\,
            I => \pulse_counter.n742\
        );

    \I__185\ : InMux
    port map (
            O => \N__2112\,
            I => \bfn_1_7_0_\
        );

    \I__184\ : InMux
    port map (
            O => \N__2109\,
            I => \pulse_counter.n728\
        );

    \I__183\ : InMux
    port map (
            O => \N__2106\,
            I => \pulse_counter.n729\
        );

    \I__182\ : InMux
    port map (
            O => \N__2103\,
            I => \pulse_counter.n730\
        );

    \I__181\ : InMux
    port map (
            O => \N__2100\,
            I => \pulse_counter.n731\
        );

    \I__180\ : InMux
    port map (
            O => \N__2097\,
            I => \pulse_counter.n732\
        );

    \I__179\ : InMux
    port map (
            O => \N__2094\,
            I => \pulse_counter.n733\
        );

    \IN_MUX_bfv_6_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_7_0_\
        );

    \IN_MUX_bfv_6_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \row_counter.n703\,
            carryinitout => \bfn_6_8_0_\
        );

    \IN_MUX_bfv_6_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \row_counter.n711\,
            carryinitout => \bfn_6_9_0_\
        );

    \IN_MUX_bfv_5_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_7_0_\
        );

    \IN_MUX_bfv_5_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \row_counter.n750\,
            carryinitout => \bfn_5_8_0_\
        );

    \IN_MUX_bfv_2_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_7_0_\
        );

    \IN_MUX_bfv_2_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pulse_counter.n719\,
            carryinitout => \bfn_2_8_0_\
        );

    \IN_MUX_bfv_2_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pulse_counter.n727\,
            carryinitout => \bfn_2_9_0_\
        );

    \IN_MUX_bfv_1_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_7_0_\
        );

    \IN_MUX_bfv_1_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pulse_counter.n735\,
            carryinitout => \bfn_1_8_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \pulse_counter.internal_count__i0_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2213\,
            in2 => \_gnd_net_\,
            in3 => \N__2112\,
            lcout => \pulse_counter.internal_count_0\,
            ltout => OPEN,
            carryin => \bfn_1_7_0_\,
            carryout => \pulse_counter.n728\,
            clk => \N__2631\,
            ce => \N__2265\,
            sr => \N__3919\
        );

    \pulse_counter.internal_count__i1_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2198\,
            in2 => \_gnd_net_\,
            in3 => \N__2109\,
            lcout => \pulse_counter.internal_count_1\,
            ltout => OPEN,
            carryin => \pulse_counter.n728\,
            carryout => \pulse_counter.n729\,
            clk => \N__2631\,
            ce => \N__2265\,
            sr => \N__3919\
        );

    \pulse_counter.internal_count__i2_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2184\,
            in2 => \_gnd_net_\,
            in3 => \N__2106\,
            lcout => \pulse_counter.internal_count_2\,
            ltout => OPEN,
            carryin => \pulse_counter.n729\,
            carryout => \pulse_counter.n730\,
            clk => \N__2631\,
            ce => \N__2265\,
            sr => \N__3919\
        );

    \pulse_counter.internal_count__i3_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2169\,
            in2 => \_gnd_net_\,
            in3 => \N__2103\,
            lcout => \pulse_counter.internal_count_3\,
            ltout => OPEN,
            carryin => \pulse_counter.n730\,
            carryout => \pulse_counter.n731\,
            clk => \N__2631\,
            ce => \N__2265\,
            sr => \N__3919\
        );

    \pulse_counter.internal_count__i4_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2154\,
            in2 => \_gnd_net_\,
            in3 => \N__2100\,
            lcout => \pulse_counter.internal_count_4\,
            ltout => OPEN,
            carryin => \pulse_counter.n731\,
            carryout => \pulse_counter.n732\,
            clk => \N__2631\,
            ce => \N__2265\,
            sr => \N__3919\
        );

    \pulse_counter.internal_count__i5_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2421\,
            in2 => \_gnd_net_\,
            in3 => \N__2097\,
            lcout => \pulse_counter.internal_count_5\,
            ltout => OPEN,
            carryin => \pulse_counter.n732\,
            carryout => \pulse_counter.n733\,
            clk => \N__2631\,
            ce => \N__2265\,
            sr => \N__3919\
        );

    \pulse_counter.internal_count__i6_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2406\,
            in2 => \_gnd_net_\,
            in3 => \N__2094\,
            lcout => \pulse_counter.internal_count_6\,
            ltout => OPEN,
            carryin => \pulse_counter.n733\,
            carryout => \pulse_counter.n734\,
            clk => \N__2631\,
            ce => \N__2265\,
            sr => \N__3919\
        );

    \pulse_counter.internal_count__i7_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2391\,
            in2 => \_gnd_net_\,
            in3 => \N__2139\,
            lcout => \pulse_counter.internal_count_7\,
            ltout => OPEN,
            carryin => \pulse_counter.n734\,
            carryout => \pulse_counter.n735\,
            clk => \N__2631\,
            ce => \N__2265\,
            sr => \N__3919\
        );

    \pulse_counter.internal_count__i8_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2376\,
            in2 => \_gnd_net_\,
            in3 => \N__2136\,
            lcout => \pulse_counter.internal_count_8\,
            ltout => OPEN,
            carryin => \bfn_1_8_0_\,
            carryout => \pulse_counter.n736\,
            clk => \N__2629\,
            ce => \N__2261\,
            sr => \N__3915\
        );

    \pulse_counter.internal_count__i9_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2361\,
            in2 => \_gnd_net_\,
            in3 => \N__2133\,
            lcout => \pulse_counter.internal_count_9\,
            ltout => OPEN,
            carryin => \pulse_counter.n736\,
            carryout => \pulse_counter.n737\,
            clk => \N__2629\,
            ce => \N__2261\,
            sr => \N__3915\
        );

    \pulse_counter.internal_count__i10_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2346\,
            in2 => \_gnd_net_\,
            in3 => \N__2130\,
            lcout => \pulse_counter.internal_count_10\,
            ltout => OPEN,
            carryin => \pulse_counter.n737\,
            carryout => \pulse_counter.n738\,
            clk => \N__2629\,
            ce => \N__2261\,
            sr => \N__3915\
        );

    \pulse_counter.internal_count__i11_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2331\,
            in2 => \_gnd_net_\,
            in3 => \N__2127\,
            lcout => \pulse_counter.internal_count_11\,
            ltout => OPEN,
            carryin => \pulse_counter.n738\,
            carryout => \pulse_counter.n739\,
            clk => \N__2629\,
            ce => \N__2261\,
            sr => \N__3915\
        );

    \pulse_counter.internal_count__i12_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2316\,
            in2 => \_gnd_net_\,
            in3 => \N__2124\,
            lcout => \pulse_counter.internal_count_12\,
            ltout => OPEN,
            carryin => \pulse_counter.n739\,
            carryout => \pulse_counter.n740\,
            clk => \N__2629\,
            ce => \N__2261\,
            sr => \N__3915\
        );

    \pulse_counter.internal_count__i13_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2301\,
            in2 => \_gnd_net_\,
            in3 => \N__2121\,
            lcout => \pulse_counter.internal_count_13\,
            ltout => OPEN,
            carryin => \pulse_counter.n740\,
            carryout => \pulse_counter.n741\,
            clk => \N__2629\,
            ce => \N__2261\,
            sr => \N__3915\
        );

    \pulse_counter.internal_count__i14_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2540\,
            in2 => \_gnd_net_\,
            in3 => \N__2118\,
            lcout => \pulse_counter.internal_count_14\,
            ltout => OPEN,
            carryin => \pulse_counter.n741\,
            carryout => \pulse_counter.n742\,
            clk => \N__2629\,
            ce => \N__2261\,
            sr => \N__3915\
        );

    \pulse_counter.internal_count__i15_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2522\,
            in2 => \_gnd_net_\,
            in3 => \N__2115\,
            lcout => \pulse_counter.internal_count_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2629\,
            ce => \N__2261\,
            sr => \N__3915\
        );

    \output_state_20_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001100010"
        )
    port map (
            in0 => \N__2243\,
            in1 => \N__2647\,
            in2 => \N__2286\,
            in3 => \N__3878\,
            lcout => output_state,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2628\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__2282\,
            in1 => \N__2646\,
            in2 => \_gnd_net_\,
            in3 => \N__3877\,
            lcout => n176,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \output_state_I_0_21_2_lut_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2244\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2232\,
            lcout => divided_pulse_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_counter.sub_8_add_2_2_lut_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__2214\,
            in1 => \N__2577\,
            in2 => \_gnd_net_\,
            in3 => \N__2202\,
            lcout => n1_adj_117,
            ltout => OPEN,
            carryin => \bfn_2_7_0_\,
            carryout => \pulse_counter.n712\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_counter.sub_8_add_2_3_lut_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__2199\,
            in1 => \N__2550\,
            in2 => \N__4218\,
            in3 => \N__2187\,
            lcout => n2_adj_99,
            ltout => OPEN,
            carryin => \pulse_counter.n712\,
            carryout => \pulse_counter.n713\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_counter.sub_8_add_2_4_lut_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__2183\,
            in1 => \N__4201\,
            in2 => \N__2613\,
            in3 => \N__2172\,
            lcout => n3_adj_118,
            ltout => OPEN,
            carryin => \pulse_counter.n713\,
            carryout => \pulse_counter.n714\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_counter.sub_8_add_2_5_lut_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__2168\,
            in1 => \N__2568\,
            in2 => \N__4219\,
            in3 => \N__2157\,
            lcout => n4_adj_116,
            ltout => OPEN,
            carryin => \pulse_counter.n714\,
            carryout => \pulse_counter.n715\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_counter.sub_8_add_2_6_lut_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__2153\,
            in1 => \N__4205\,
            in2 => \N__2739\,
            in3 => \N__2142\,
            lcout => n5_adj_120,
            ltout => OPEN,
            carryin => \pulse_counter.n715\,
            carryout => \pulse_counter.n716\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_counter.sub_8_add_2_7_lut_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__2420\,
            in1 => \N__2727\,
            in2 => \N__4220\,
            in3 => \N__2409\,
            lcout => n6_adj_119,
            ltout => OPEN,
            carryin => \pulse_counter.n716\,
            carryout => \pulse_counter.n717\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_counter.sub_8_add_2_8_lut_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__2405\,
            in1 => \N__2757\,
            in2 => \N__4212\,
            in3 => \N__2394\,
            lcout => n7,
            ltout => OPEN,
            carryin => \pulse_counter.n717\,
            carryout => \pulse_counter.n718\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_counter.sub_8_add_2_9_lut_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__2390\,
            in1 => \N__2706\,
            in2 => \N__4221\,
            in3 => \N__2379\,
            lcout => n8,
            ltout => OPEN,
            carryin => \pulse_counter.n718\,
            carryout => \pulse_counter.n719\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_counter.sub_8_add_2_10_lut_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__2375\,
            in1 => \N__2718\,
            in2 => \N__4213\,
            in3 => \N__2364\,
            lcout => n9,
            ltout => OPEN,
            carryin => \bfn_2_8_0_\,
            carryout => \pulse_counter.n720\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_counter.sub_8_add_2_11_lut_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__2360\,
            in1 => \N__2748\,
            in2 => \N__4216\,
            in3 => \N__2349\,
            lcout => n10,
            ltout => OPEN,
            carryin => \pulse_counter.n720\,
            carryout => \pulse_counter.n721\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_counter.sub_8_add_2_12_lut_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__2345\,
            in1 => \N__2766\,
            in2 => \N__4214\,
            in3 => \N__2334\,
            lcout => n11,
            ltout => OPEN,
            carryin => \pulse_counter.n721\,
            carryout => \pulse_counter.n722\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_counter.sub_8_add_2_13_lut_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__2330\,
            in1 => \N__2427\,
            in2 => \N__4217\,
            in3 => \N__2319\,
            lcout => n12,
            ltout => OPEN,
            carryin => \pulse_counter.n722\,
            carryout => \pulse_counter.n723\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_counter.sub_8_add_2_14_lut_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__2315\,
            in1 => \N__2559\,
            in2 => \N__4215\,
            in3 => \N__2304\,
            lcout => \pulse_counter.n13\,
            ltout => OPEN,
            carryin => \pulse_counter.n723\,
            carryout => \pulse_counter.n724\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_counter.sub_8_add_2_15_lut_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__2300\,
            in1 => \N__4189\,
            in2 => \N__2658\,
            in3 => \N__2289\,
            lcout => n14,
            ltout => OPEN,
            carryin => \pulse_counter.n724\,
            carryout => \pulse_counter.n725\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_counter.sub_8_add_2_16_lut_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__2541\,
            in1 => \N__4197\,
            in2 => \N__2601\,
            in3 => \N__2526\,
            lcout => n15,
            ltout => OPEN,
            carryin => \pulse_counter.n725\,
            carryout => \pulse_counter.n726\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_counter.sub_8_add_2_17_lut_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__2523\,
            in1 => \N__4190\,
            in2 => \N__2589\,
            in3 => \N__2508\,
            lcout => n16,
            ltout => OPEN,
            carryin => \pulse_counter.n726\,
            carryout => \pulse_counter.n727\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_counter.sub_8_add_2_18_lut_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110111011110"
        )
    port map (
            in0 => \N__4119\,
            in1 => \N__2505\,
            in2 => \_gnd_net_\,
            in3 => \N__2499\,
            lcout => n787,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i732_2_lut_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2496\,
            in2 => \_gnd_net_\,
            in3 => \N__2487\,
            lcout => OPEN,
            ltout => \n795_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i754_4_lut_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__2478\,
            in1 => \N__2469\,
            in2 => \N__2463\,
            in3 => \N__2460\,
            lcout => OPEN,
            ltout => \n817_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i762_4_lut_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__2451\,
            in1 => \N__2445\,
            in2 => \N__2439\,
            in3 => \N__2436\,
            lcout => OPEN,
            ltout => \n825_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pulse_counter.internal_count_reached_18_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101011"
        )
    port map (
            in0 => \N__2649\,
            in1 => \N__2883\,
            in2 => \N__2430\,
            in3 => \N__3879\,
            lcout => count_done,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2630\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.output_enable_I_0_i12_2_lut_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2781\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4622\,
            lcout => sr_divider_data_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.output_enable_I_0_i14_2_lut_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4623\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3027\,
            lcout => sr_divider_data_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_signal_19_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__3880\,
            in1 => \N__2648\,
            in2 => \_gnd_net_\,
            in3 => \N__3828\,
            lcout => reset_signal,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2630\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.output_enable_I_0_i3_2_lut_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4591\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3350\,
            lcout => sr_divider_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.output_enable_I_0_i15_2_lut_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4587\,
            in2 => \_gnd_net_\,
            in3 => \N__2808\,
            lcout => sr_divider_data_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.output_enable_I_0_i16_2_lut_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4588\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2793\,
            lcout => sr_divider_data_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.output_enable_I_0_i1_2_lut_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4589\,
            in2 => \_gnd_net_\,
            in3 => \N__3393\,
            lcout => sr_divider_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.output_enable_I_0_i4_2_lut_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4592\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3165\,
            lcout => sr_divider_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.output_enable_I_0_i13_2_lut_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3047\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4586\,
            lcout => sr_divider_data_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.output_enable_I_0_i2_2_lut_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__4590\,
            in1 => \N__3375\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => sr_divider_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.output_enable_I_0_i11_2_lut_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4585\,
            in2 => \_gnd_net_\,
            in3 => \N__2976\,
            lcout => sr_divider_data_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.output_enable_I_0_i7_2_lut_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__2943\,
            in1 => \N__4548\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => sr_divider_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.output_enable_I_0_i10_2_lut_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4545\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2996\,
            lcout => sr_divider_data_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.output_enable_I_0_i5_2_lut_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3140\,
            in2 => \_gnd_net_\,
            in3 => \N__4546\,
            lcout => sr_divider_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.output_enable_I_0_i6_2_lut_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4547\,
            in2 => \_gnd_net_\,
            in3 => \N__2958\,
            lcout => sr_divider_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.output_enable_I_0_i9_2_lut_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4550\,
            in2 => \_gnd_net_\,
            in3 => \N__3012\,
            lcout => sr_divider_data_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.output_enable_I_0_i8_2_lut_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4549\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2927\,
            lcout => sr_divider_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i718_2_lut_LC_3_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2697\,
            in2 => \_gnd_net_\,
            in3 => \N__2691\,
            lcout => n781,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i760_4_lut_LC_3_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__2685\,
            in1 => \N__2679\,
            in2 => \N__2673\,
            in3 => \N__2664\,
            lcout => OPEN,
            ltout => \n823_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i764_4_lut_LC_3_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__2904\,
            in1 => \N__2898\,
            in2 => \N__2892\,
            in3 => \N__2889\,
            lcout => n827,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i355_2_lut_3_lut_LC_3_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__3892\,
            in1 => \N__2877\,
            in2 => \_gnd_net_\,
            in3 => \N__2836\,
            lcout => n345,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_5_LC_3_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__3891\,
            in1 => \N__2876\,
            in2 => \_gnd_net_\,
            in3 => \N__2835\,
            lcout => n171,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.shifted_data_i11_LC_3_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__3289\,
            in1 => \N__2779\,
            in2 => \N__3236\,
            in3 => \N__2975\,
            lcout => shifted_data_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4708\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__2855\,
            in1 => \N__2837\,
            in2 => \_gnd_net_\,
            in3 => \N__3893\,
            lcout => n169,
            ltout => \n169_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.shifted_data_i14_LC_3_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__3294\,
            in1 => \N__2806\,
            in2 => \N__2859\,
            in3 => \N__3026\,
            lcout => shifted_data_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4708\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i340_2_lut_3_lut_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__2856\,
            in1 => \N__2838\,
            in2 => \_gnd_net_\,
            in3 => \N__3894\,
            lcout => n330,
            ltout => \n330_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.shifted_data_i15_LC_3_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__3211\,
            in1 => \N__2792\,
            in2 => \N__2811\,
            in3 => \N__2807\,
            lcout => shifted_data_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4708\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.shifted_data_i12_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__2780\,
            in1 => \N__3290\,
            in2 => \N__3048\,
            in3 => \N__3210\,
            lcout => shifted_data_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4708\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.shifted_data_i13_LC_3_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__3043\,
            in1 => \N__3212\,
            in2 => \N__3315\,
            in3 => \N__3025\,
            lcout => shifted_data_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4708\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.shifted_data_i8_LC_3_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__2923\,
            in1 => \N__3221\,
            in2 => \N__3316\,
            in3 => \N__3010\,
            lcout => shifted_data_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4709\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.shifted_data_i6_LC_3_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__2956\,
            in1 => \N__3297\,
            in2 => \N__3238\,
            in3 => \N__2941\,
            lcout => shifted_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4709\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.shifted_data_i9_LC_3_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__3302\,
            in1 => \N__3222\,
            in2 => \N__2997\,
            in3 => \N__3011\,
            lcout => shifted_data_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4709\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.shifted_data_i10_LC_3_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__2992\,
            in1 => \N__3295\,
            in2 => \N__3237\,
            in3 => \N__2974\,
            lcout => shifted_data_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4709\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.shifted_data_i5_LC_3_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__3296\,
            in1 => \N__3216\,
            in2 => \N__3141\,
            in3 => \N__2957\,
            lcout => shifted_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4709\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.shifted_data_i7_LC_3_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__3220\,
            in1 => \N__2942\,
            in2 => \N__2928\,
            in3 => \N__3298\,
            lcout => shifted_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4709\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.shifted_data_i0_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__3416\,
            in1 => \N__4964\,
            in2 => \N__4878\,
            in3 => \N__3109\,
            lcout => shifted_data_0_adj_115,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4716\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_counter.internal_count__i0_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3620\,
            in2 => \_gnd_net_\,
            in3 => \N__2907\,
            lcout => \row_counter.internal_count_0\,
            ltout => OPEN,
            carryin => \bfn_5_7_0_\,
            carryout => \row_counter.n743\,
            clk => \N__3803\,
            ce => \N__3438\,
            sr => \N__3924\
        );

    \row_counter.internal_count__i1_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3596\,
            in2 => \_gnd_net_\,
            in3 => \N__3075\,
            lcout => \row_counter.internal_count_1\,
            ltout => OPEN,
            carryin => \row_counter.n743\,
            carryout => \row_counter.n744\,
            clk => \N__3803\,
            ce => \N__3438\,
            sr => \N__3924\
        );

    \row_counter.internal_count__i2_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3573\,
            in2 => \_gnd_net_\,
            in3 => \N__3072\,
            lcout => \row_counter.internal_count_2\,
            ltout => OPEN,
            carryin => \row_counter.n744\,
            carryout => \row_counter.n745\,
            clk => \N__3803\,
            ce => \N__3438\,
            sr => \N__3924\
        );

    \row_counter.internal_count__i3_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3551\,
            in2 => \_gnd_net_\,
            in3 => \N__3069\,
            lcout => \row_counter.internal_count_3\,
            ltout => OPEN,
            carryin => \row_counter.n745\,
            carryout => \row_counter.n746\,
            clk => \N__3803\,
            ce => \N__3438\,
            sr => \N__3924\
        );

    \row_counter.internal_count__i4_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3537\,
            in2 => \_gnd_net_\,
            in3 => \N__3066\,
            lcout => \row_counter.internal_count_4\,
            ltout => OPEN,
            carryin => \row_counter.n746\,
            carryout => \row_counter.n747\,
            clk => \N__3803\,
            ce => \N__3438\,
            sr => \N__3924\
        );

    \row_counter.internal_count__i5_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3512\,
            in2 => \_gnd_net_\,
            in3 => \N__3063\,
            lcout => \row_counter.internal_count_5\,
            ltout => OPEN,
            carryin => \row_counter.n747\,
            carryout => \row_counter.n748\,
            clk => \N__3803\,
            ce => \N__3438\,
            sr => \N__3924\
        );

    \row_counter.internal_count__i6_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3498\,
            in2 => \_gnd_net_\,
            in3 => \N__3060\,
            lcout => \row_counter.internal_count_6\,
            ltout => OPEN,
            carryin => \row_counter.n748\,
            carryout => \row_counter.n749\,
            clk => \N__3803\,
            ce => \N__3438\,
            sr => \N__3924\
        );

    \row_counter.internal_count__i7_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3483\,
            in2 => \_gnd_net_\,
            in3 => \N__3057\,
            lcout => \row_counter.internal_count_7\,
            ltout => OPEN,
            carryin => \row_counter.n749\,
            carryout => \row_counter.n750\,
            clk => \N__3803\,
            ce => \N__3438\,
            sr => \N__3924\
        );

    \row_counter.internal_count__i8_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3756\,
            in2 => \_gnd_net_\,
            in3 => \N__3054\,
            lcout => \row_counter.internal_count_8\,
            ltout => OPEN,
            carryin => \bfn_5_8_0_\,
            carryout => \row_counter.n751\,
            clk => \N__3802\,
            ce => \N__3437\,
            sr => \N__3923\
        );

    \row_counter.internal_count__i9_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3740\,
            in2 => \_gnd_net_\,
            in3 => \N__3051\,
            lcout => \row_counter.internal_count_9\,
            ltout => OPEN,
            carryin => \row_counter.n751\,
            carryout => \row_counter.n752\,
            clk => \N__3802\,
            ce => \N__3437\,
            sr => \N__3923\
        );

    \row_counter.internal_count__i10_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3723\,
            in2 => \_gnd_net_\,
            in3 => \N__3093\,
            lcout => \row_counter.internal_count_10\,
            ltout => OPEN,
            carryin => \row_counter.n752\,
            carryout => \row_counter.n753\,
            clk => \N__3802\,
            ce => \N__3437\,
            sr => \N__3923\
        );

    \row_counter.internal_count__i11_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3708\,
            in2 => \_gnd_net_\,
            in3 => \N__3090\,
            lcout => \row_counter.internal_count_11\,
            ltout => OPEN,
            carryin => \row_counter.n753\,
            carryout => \row_counter.n754\,
            clk => \N__3802\,
            ce => \N__3437\,
            sr => \N__3923\
        );

    \row_counter.internal_count__i12_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3693\,
            in2 => \_gnd_net_\,
            in3 => \N__3087\,
            lcout => \row_counter.internal_count_12\,
            ltout => OPEN,
            carryin => \row_counter.n754\,
            carryout => \row_counter.n755\,
            clk => \N__3802\,
            ce => \N__3437\,
            sr => \N__3923\
        );

    \row_counter.internal_count__i13_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3678\,
            in2 => \_gnd_net_\,
            in3 => \N__3084\,
            lcout => \row_counter.internal_count_13\,
            ltout => OPEN,
            carryin => \row_counter.n755\,
            carryout => \row_counter.n756\,
            clk => \N__3802\,
            ce => \N__3437\,
            sr => \N__3923\
        );

    \row_counter.internal_count__i14_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3663\,
            in2 => \_gnd_net_\,
            in3 => \N__3081\,
            lcout => \row_counter.internal_count_14\,
            ltout => OPEN,
            carryin => \row_counter.n756\,
            carryout => \row_counter.n757\,
            clk => \N__3802\,
            ce => \N__3437\,
            sr => \N__3923\
        );

    \row_counter.internal_count__i15_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3648\,
            in2 => \_gnd_net_\,
            in3 => \N__3078\,
            lcout => \row_counter.internal_count_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3802\,
            ce => \N__3437\,
            sr => \N__3923\
        );

    \CONSTANT_ONE_LUT4_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.output_enable_I_0_i1_2_lut_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3114\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4619\,
            lcout => sr_row_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.output_enable_I_0_i5_2_lut_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4620\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4416\,
            lcout => sr_row_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.output_enable_I_0_i8_2_lut_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4621\,
            in2 => \_gnd_net_\,
            in3 => \N__4320\,
            lcout => sr_row_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_7_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__3456\,
            in1 => \N__3820\,
            in2 => \_gnd_net_\,
            in3 => \N__3913\,
            lcout => n189,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.shifted_data_i1_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__3389\,
            in1 => \N__3318\,
            in2 => \N__3374\,
            in3 => \N__3242\,
            lcout => shifted_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.shifted_data_i0_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__3317\,
            in1 => \N__3420\,
            in2 => \N__3248\,
            in3 => \N__3388\,
            lcout => shifted_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.shifted_data_i3_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__3244\,
            in1 => \N__3343\,
            in2 => \N__3164\,
            in3 => \N__3320\,
            lcout => shifted_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.shifted_data_i2_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__3243\,
            in1 => \N__3367\,
            in2 => \N__3351\,
            in3 => \N__3319\,
            lcout => shifted_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \divider_sr.shifted_data_i4_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__3324\,
            in1 => \N__3133\,
            in2 => \N__3252\,
            in3 => \N__3160\,
            lcout => shifted_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4712\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.shifted_data_i1_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__4965\,
            in1 => \N__3631\,
            in2 => \N__4879\,
            in3 => \N__3110\,
            lcout => shifted_data_1_adj_114,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4717\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.output_enable_I_0_i2_2_lut_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3633\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4645\,
            lcout => sr_row_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.shifted_data_i2_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__4966\,
            in1 => \N__4450\,
            in2 => \N__4880\,
            in3 => \N__3632\,
            lcout => shifted_data_2_adj_113,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4717\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_counter.sub_8_add_2_2_lut_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__3621\,
            in1 => \N__3609\,
            in2 => \_gnd_net_\,
            in3 => \N__3600\,
            lcout => n1,
            ltout => OPEN,
            carryin => \bfn_6_7_0_\,
            carryout => \row_counter.n696\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_counter.sub_8_add_2_3_lut_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__3597\,
            in1 => \N__4120\,
            in2 => \N__3585\,
            in3 => \N__3576\,
            lcout => n2,
            ltout => OPEN,
            carryin => \row_counter.n696\,
            carryout => \row_counter.n697\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_counter.sub_8_add_2_4_lut_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__3572\,
            in1 => \N__4434\,
            in2 => \N__4143\,
            in3 => \N__3558\,
            lcout => n3,
            ltout => OPEN,
            carryin => \row_counter.n697\,
            carryout => \row_counter.n698\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_counter.sub_8_add_2_5_lut_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__3555\,
            in1 => \N__4124\,
            in2 => \N__4464\,
            in3 => \N__3540\,
            lcout => n4,
            ltout => OPEN,
            carryin => \row_counter.n698\,
            carryout => \row_counter.n699\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_counter.sub_8_add_2_6_lut_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__3536\,
            in1 => \N__3525\,
            in2 => \N__4144\,
            in3 => \N__3516\,
            lcout => n5,
            ltout => OPEN,
            carryin => \row_counter.n699\,
            carryout => \row_counter.n700\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_counter.sub_8_add_2_7_lut_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__3513\,
            in1 => \N__4128\,
            in2 => \N__4662\,
            in3 => \N__3501\,
            lcout => n6,
            ltout => OPEN,
            carryin => \row_counter.n700\,
            carryout => \row_counter.n701\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_counter.sub_8_add_2_8_lut_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__3497\,
            in1 => \N__4008\,
            in2 => \N__4145\,
            in3 => \N__3486\,
            lcout => n7_adj_121,
            ltout => OPEN,
            carryin => \row_counter.n701\,
            carryout => \row_counter.n702\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_counter.sub_8_add_2_9_lut_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__3482\,
            in1 => \N__4132\,
            in2 => \N__3471\,
            in3 => \N__3459\,
            lcout => n8_adj_122,
            ltout => OPEN,
            carryin => \row_counter.n702\,
            carryout => \row_counter.n703\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_counter.sub_8_add_2_10_lut_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__3755\,
            in1 => \N__4014\,
            in2 => \N__4111\,
            in3 => \N__3744\,
            lcout => n9_adj_123,
            ltout => OPEN,
            carryin => \bfn_6_8_0_\,
            carryout => \row_counter.n704\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_counter.sub_8_add_2_11_lut_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__3741\,
            in1 => \N__3999\,
            in2 => \N__4115\,
            in3 => \N__3726\,
            lcout => n10_adj_124,
            ltout => OPEN,
            carryin => \row_counter.n704\,
            carryout => \row_counter.n705\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_counter.sub_8_add_2_12_lut_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__3722\,
            in1 => \N__4236\,
            in2 => \N__4112\,
            in3 => \N__3711\,
            lcout => n11_adj_125,
            ltout => OPEN,
            carryin => \row_counter.n705\,
            carryout => \row_counter.n706\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_counter.sub_8_add_2_13_lut_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__3707\,
            in1 => \N__4287\,
            in2 => \N__4116\,
            in3 => \N__3696\,
            lcout => n12_adj_126,
            ltout => OPEN,
            carryin => \row_counter.n706\,
            carryout => \row_counter.n707\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_counter.sub_8_add_2_14_lut_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__3692\,
            in1 => \N__5034\,
            in2 => \N__4113\,
            in3 => \N__3681\,
            lcout => \row_counter.n13\,
            ltout => OPEN,
            carryin => \row_counter.n707\,
            carryout => \row_counter.n708\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_counter.sub_8_add_2_15_lut_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__3677\,
            in1 => \N__4269\,
            in2 => \N__4117\,
            in3 => \N__3666\,
            lcout => n14_adj_127,
            ltout => OPEN,
            carryin => \row_counter.n708\,
            carryout => \row_counter.n709\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_counter.sub_8_add_2_16_lut_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__3662\,
            in1 => \N__4296\,
            in2 => \N__4114\,
            in3 => \N__3651\,
            lcout => n15_adj_128,
            ltout => OPEN,
            carryin => \row_counter.n709\,
            carryout => \row_counter.n710\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_counter.sub_8_add_2_17_lut_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__3647\,
            in1 => \N__4278\,
            in2 => \N__4118\,
            in3 => \N__3636\,
            lcout => n16_adj_129,
            ltout => OPEN,
            carryin => \row_counter.n710\,
            carryout => \row_counter.n711\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_counter.sub_8_add_2_18_lut_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__4227\,
            in1 => \N__4062\,
            in2 => \_gnd_net_\,
            in3 => \N__4017\,
            lcout => n775,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.output_enable_I_0_i9_2_lut_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4648\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5049\,
            lcout => sr_row_data_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.output_enable_I_0_i7_2_lut_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4647\,
            in2 => \_gnd_net_\,
            in3 => \N__4341\,
            lcout => sr_row_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.output_enable_I_0_i10_2_lut_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4646\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4754\,
            lcout => sr_row_data_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i748_2_lut_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3993\,
            in2 => \_gnd_net_\,
            in3 => \N__3984\,
            lcout => OPEN,
            ltout => \n811_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i768_4_lut_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3975\,
            in1 => \N__3966\,
            in2 => \N__3960\,
            in3 => \N__3957\,
            lcout => OPEN,
            ltout => \n831_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i772_4_lut_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3948\,
            in1 => \N__3939\,
            in2 => \N__3933\,
            in3 => \N__3930\,
            lcout => OPEN,
            ltout => \n835_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_counter.internal_count_reached_18_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000100011"
        )
    port map (
            in0 => \N__3821\,
            in1 => \N__3914\,
            in2 => \N__3831\,
            in3 => \N__4347\,
            lcout => row_complete,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3804\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.output_enable_I_0_i15_2_lut_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4630\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4248\,
            lcout => sr_row_data_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.output_enable_I_0_i12_2_lut_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5003\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4628\,
            lcout => sr_row_data_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.shifted_data_i11_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__4961\,
            in1 => \N__5002\,
            in2 => \N__4862\,
            in3 => \N__4733\,
            lcout => shifted_data_11_adj_104,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4711\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.output_enable_I_0_i16_2_lut_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__4259\,
            in1 => \N__4631\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => sr_row_data_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.output_enable_I_0_i14_2_lut_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4629\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5024\,
            lcout => sr_row_data_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.shifted_data_i15_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__4247\,
            in1 => \N__4963\,
            in2 => \N__4260\,
            in3 => \N__4835\,
            lcout => shifted_data_15_adj_100,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4711\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.shifted_data_i14_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__4962\,
            in1 => \N__4246\,
            in2 => \N__4863\,
            in3 => \N__5023\,
            lcout => shifted_data_14_adj_101,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4711\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.output_enable_I_0_i11_2_lut_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4734\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4627\,
            lcout => sr_row_data_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.shifted_data_i3_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__4976\,
            in1 => \N__4480\,
            in2 => \N__4877\,
            in3 => \N__4451\,
            lcout => shifted_data_3_adj_112,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4719\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.shifted_data_i5_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__4408\,
            in1 => \N__4872\,
            in2 => \N__4977\,
            in3 => \N__4675\,
            lcout => shifted_data_5_adj_110,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4718\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.output_enable_I_0_i3_2_lut_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4650\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4452\,
            lcout => sr_row_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i740_2_lut_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4428\,
            in2 => \_gnd_net_\,
            in3 => \N__4422\,
            lcout => n803,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.shifted_data_i6_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__4676\,
            in1 => \N__4975\,
            in2 => \N__4881\,
            in3 => \N__4336\,
            lcout => shifted_data_6_adj_109,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4718\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.shifted_data_i4_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__4871\,
            in1 => \N__4971\,
            in2 => \N__4488\,
            in3 => \N__4409\,
            lcout => shifted_data_4_adj_111,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4718\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i730_4_lut_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4395\,
            in1 => \N__4389\,
            in2 => \N__4383\,
            in3 => \N__4374\,
            lcout => OPEN,
            ltout => \n793_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i766_4_lut_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4368\,
            in1 => \N__4362\,
            in2 => \N__4356\,
            in3 => \N__4353\,
            lcout => n829,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.shifted_data_i7_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__4970\,
            in1 => \N__4312\,
            in2 => \N__4876\,
            in3 => \N__4337\,
            lcout => shifted_data_7_adj_108,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4715\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.shifted_data_i8_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__4924\,
            in1 => \N__5047\,
            in2 => \N__4828\,
            in3 => \N__4313\,
            lcout => shifted_data_8_adj_107,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4714\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.shifted_data_i9_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__5048\,
            in1 => \N__4798\,
            in2 => \N__4755\,
            in3 => \N__4925\,
            lcout => shifted_data_9_adj_106,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4714\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.output_enable_I_0_i13_2_lut_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4649\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4989\,
            lcout => sr_row_data_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.shifted_data_i13_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__4840\,
            in1 => \N__4988\,
            in2 => \N__5025\,
            in3 => \N__4969\,
            lcout => shifted_data_13_adj_102,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4713\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.shifted_data_i12_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__4839\,
            in1 => \N__4987\,
            in2 => \N__5007\,
            in3 => \N__4968\,
            lcout => shifted_data_12_adj_103,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4713\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.shifted_data_i10_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__4967\,
            in1 => \N__4732\,
            in2 => \N__4864\,
            in3 => \N__4753\,
            lcout => shifted_data_10_adj_105,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4713\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.output_enable_I_0_i6_2_lut_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4677\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4544\,
            lcout => sr_row_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_sr.output_enable_I_0_i4_2_lut_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4543\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4484\,
            lcout => sr_row_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
