// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Aug 2 2023 08:20:12

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    sr_sel_row,
    sr_sel_div,
    sr_clk,
    row_completed,
    en_internals,
    divide_enable,
    sr_reset,
    laser_pulse,
    sr_data,
    en_rowpack,
    divided_pulse,
    constant_v);

    input sr_sel_row;
    input sr_sel_div;
    input sr_clk;
    output row_completed;
    input en_internals;
    input divide_enable;
    input sr_reset;
    input laser_pulse;
    input sr_data;
    input en_rowpack;
    output divided_pulse;
    input constant_v;

    wire N__5170;
    wire N__5169;
    wire N__5168;
    wire N__5160;
    wire N__5159;
    wire N__5158;
    wire N__5149;
    wire N__5148;
    wire N__5147;
    wire N__5140;
    wire N__5139;
    wire N__5138;
    wire N__5131;
    wire N__5130;
    wire N__5129;
    wire N__5122;
    wire N__5121;
    wire N__5120;
    wire N__5113;
    wire N__5112;
    wire N__5111;
    wire N__5104;
    wire N__5103;
    wire N__5102;
    wire N__5095;
    wire N__5094;
    wire N__5093;
    wire N__5086;
    wire N__5085;
    wire N__5084;
    wire N__5077;
    wire N__5076;
    wire N__5075;
    wire N__5068;
    wire N__5067;
    wire N__5066;
    wire N__5049;
    wire N__5048;
    wire N__5047;
    wire N__5044;
    wire N__5039;
    wire N__5034;
    wire N__5031;
    wire N__5028;
    wire N__5025;
    wire N__5024;
    wire N__5023;
    wire N__5020;
    wire N__5015;
    wire N__5012;
    wire N__5007;
    wire N__5004;
    wire N__5003;
    wire N__5002;
    wire N__4999;
    wire N__4994;
    wire N__4989;
    wire N__4988;
    wire N__4987;
    wire N__4980;
    wire N__4977;
    wire N__4976;
    wire N__4975;
    wire N__4972;
    wire N__4971;
    wire N__4970;
    wire N__4969;
    wire N__4968;
    wire N__4967;
    wire N__4966;
    wire N__4965;
    wire N__4964;
    wire N__4963;
    wire N__4962;
    wire N__4961;
    wire N__4958;
    wire N__4951;
    wire N__4948;
    wire N__4941;
    wire N__4936;
    wire N__4933;
    wire N__4926;
    wire N__4925;
    wire N__4924;
    wire N__4917;
    wire N__4914;
    wire N__4909;
    wire N__4906;
    wire N__4901;
    wire N__4896;
    wire N__4891;
    wire N__4888;
    wire N__4881;
    wire N__4880;
    wire N__4879;
    wire N__4878;
    wire N__4877;
    wire N__4876;
    wire N__4873;
    wire N__4872;
    wire N__4871;
    wire N__4868;
    wire N__4865;
    wire N__4864;
    wire N__4863;
    wire N__4862;
    wire N__4859;
    wire N__4856;
    wire N__4853;
    wire N__4846;
    wire N__4841;
    wire N__4840;
    wire N__4839;
    wire N__4836;
    wire N__4835;
    wire N__4832;
    wire N__4829;
    wire N__4828;
    wire N__4825;
    wire N__4822;
    wire N__4819;
    wire N__4814;
    wire N__4809;
    wire N__4806;
    wire N__4799;
    wire N__4798;
    wire N__4795;
    wire N__4792;
    wire N__4787;
    wire N__4778;
    wire N__4773;
    wire N__4770;
    wire N__4765;
    wire N__4762;
    wire N__4755;
    wire N__4754;
    wire N__4753;
    wire N__4750;
    wire N__4747;
    wire N__4744;
    wire N__4741;
    wire N__4734;
    wire N__4733;
    wire N__4732;
    wire N__4727;
    wire N__4724;
    wire N__4719;
    wire N__4718;
    wire N__4717;
    wire N__4716;
    wire N__4715;
    wire N__4714;
    wire N__4713;
    wire N__4712;
    wire N__4711;
    wire N__4710;
    wire N__4709;
    wire N__4708;
    wire N__4683;
    wire N__4680;
    wire N__4677;
    wire N__4676;
    wire N__4675;
    wire N__4672;
    wire N__4667;
    wire N__4662;
    wire N__4659;
    wire N__4656;
    wire N__4653;
    wire N__4650;
    wire N__4649;
    wire N__4648;
    wire N__4647;
    wire N__4646;
    wire N__4645;
    wire N__4642;
    wire N__4639;
    wire N__4632;
    wire N__4631;
    wire N__4630;
    wire N__4629;
    wire N__4628;
    wire N__4627;
    wire N__4624;
    wire N__4623;
    wire N__4622;
    wire N__4621;
    wire N__4620;
    wire N__4619;
    wire N__4612;
    wire N__4601;
    wire N__4598;
    wire N__4593;
    wire N__4592;
    wire N__4591;
    wire N__4590;
    wire N__4589;
    wire N__4588;
    wire N__4587;
    wire N__4586;
    wire N__4585;
    wire N__4578;
    wire N__4573;
    wire N__4568;
    wire N__4551;
    wire N__4550;
    wire N__4549;
    wire N__4548;
    wire N__4547;
    wire N__4546;
    wire N__4545;
    wire N__4544;
    wire N__4543;
    wire N__4540;
    wire N__4533;
    wire N__4520;
    wire N__4515;
    wire N__4512;
    wire N__4507;
    wire N__4504;
    wire N__4501;
    wire N__4498;
    wire N__4491;
    wire N__4488;
    wire N__4485;
    wire N__4484;
    wire N__4481;
    wire N__4480;
    wire N__4477;
    wire N__4474;
    wire N__4471;
    wire N__4464;
    wire N__4461;
    wire N__4458;
    wire N__4455;
    wire N__4452;
    wire N__4451;
    wire N__4450;
    wire N__4447;
    wire N__4444;
    wire N__4441;
    wire N__4434;
    wire N__4431;
    wire N__4428;
    wire N__4425;
    wire N__4422;
    wire N__4419;
    wire N__4416;
    wire N__4413;
    wire N__4410;
    wire N__4409;
    wire N__4408;
    wire N__4405;
    wire N__4400;
    wire N__4395;
    wire N__4392;
    wire N__4389;
    wire N__4386;
    wire N__4383;
    wire N__4380;
    wire N__4377;
    wire N__4374;
    wire N__4371;
    wire N__4368;
    wire N__4365;
    wire N__4362;
    wire N__4359;
    wire N__4356;
    wire N__4353;
    wire N__4350;
    wire N__4347;
    wire N__4344;
    wire N__4341;
    wire N__4338;
    wire N__4337;
    wire N__4336;
    wire N__4333;
    wire N__4330;
    wire N__4327;
    wire N__4320;
    wire N__4317;
    wire N__4314;
    wire N__4313;
    wire N__4312;
    wire N__4309;
    wire N__4306;
    wire N__4303;
    wire N__4296;
    wire N__4293;
    wire N__4290;
    wire N__4287;
    wire N__4284;
    wire N__4281;
    wire N__4278;
    wire N__4275;
    wire N__4272;
    wire N__4269;
    wire N__4266;
    wire N__4263;
    wire N__4260;
    wire N__4259;
    wire N__4256;
    wire N__4251;
    wire N__4248;
    wire N__4247;
    wire N__4246;
    wire N__4239;
    wire N__4236;
    wire N__4233;
    wire N__4230;
    wire N__4227;
    wire N__4224;
    wire N__4221;
    wire N__4220;
    wire N__4219;
    wire N__4218;
    wire N__4217;
    wire N__4216;
    wire N__4215;
    wire N__4214;
    wire N__4213;
    wire N__4212;
    wire N__4209;
    wire N__4206;
    wire N__4205;
    wire N__4202;
    wire N__4201;
    wire N__4198;
    wire N__4197;
    wire N__4194;
    wire N__4191;
    wire N__4190;
    wire N__4189;
    wire N__4186;
    wire N__4183;
    wire N__4180;
    wire N__4177;
    wire N__4164;
    wire N__4157;
    wire N__4146;
    wire N__4145;
    wire N__4144;
    wire N__4143;
    wire N__4140;
    wire N__4133;
    wire N__4132;
    wire N__4129;
    wire N__4128;
    wire N__4125;
    wire N__4124;
    wire N__4121;
    wire N__4120;
    wire N__4119;
    wire N__4118;
    wire N__4117;
    wire N__4116;
    wire N__4115;
    wire N__4114;
    wire N__4113;
    wire N__4112;
    wire N__4111;
    wire N__4108;
    wire N__4105;
    wire N__4090;
    wire N__4087;
    wire N__4084;
    wire N__4081;
    wire N__4078;
    wire N__4075;
    wire N__4072;
    wire N__4069;
    wire N__4066;
    wire N__4063;
    wire N__4062;
    wire N__4059;
    wire N__4054;
    wire N__4051;
    wire N__4042;
    wire N__4033;
    wire N__4030;
    wire N__4017;
    wire N__4014;
    wire N__4011;
    wire N__4008;
    wire N__4005;
    wire N__4002;
    wire N__3999;
    wire N__3996;
    wire N__3993;
    wire N__3990;
    wire N__3987;
    wire N__3984;
    wire N__3981;
    wire N__3978;
    wire N__3975;
    wire N__3972;
    wire N__3969;
    wire N__3966;
    wire N__3963;
    wire N__3960;
    wire N__3957;
    wire N__3954;
    wire N__3951;
    wire N__3948;
    wire N__3945;
    wire N__3942;
    wire N__3939;
    wire N__3936;
    wire N__3933;
    wire N__3930;
    wire N__3927;
    wire N__3924;
    wire N__3923;
    wire N__3920;
    wire N__3919;
    wire N__3916;
    wire N__3915;
    wire N__3914;
    wire N__3913;
    wire N__3910;
    wire N__3907;
    wire N__3904;
    wire N__3901;
    wire N__3898;
    wire N__3895;
    wire N__3894;
    wire N__3893;
    wire N__3892;
    wire N__3891;
    wire N__3886;
    wire N__3881;
    wire N__3880;
    wire N__3879;
    wire N__3878;
    wire N__3877;
    wire N__3872;
    wire N__3867;
    wire N__3862;
    wire N__3859;
    wire N__3856;
    wire N__3851;
    wire N__3846;
    wire N__3831;
    wire N__3828;
    wire N__3825;
    wire N__3822;
    wire N__3821;
    wire N__3820;
    wire N__3817;
    wire N__3814;
    wire N__3811;
    wire N__3804;
    wire N__3803;
    wire N__3802;
    wire N__3799;
    wire N__3796;
    wire N__3793;
    wire N__3790;
    wire N__3789;
    wire N__3786;
    wire N__3783;
    wire N__3780;
    wire N__3777;
    wire N__3774;
    wire N__3771;
    wire N__3768;
    wire N__3765;
    wire N__3756;
    wire N__3755;
    wire N__3752;
    wire N__3749;
    wire N__3744;
    wire N__3741;
    wire N__3740;
    wire N__3737;
    wire N__3734;
    wire N__3731;
    wire N__3726;
    wire N__3723;
    wire N__3722;
    wire N__3719;
    wire N__3716;
    wire N__3711;
    wire N__3708;
    wire N__3707;
    wire N__3704;
    wire N__3701;
    wire N__3696;
    wire N__3693;
    wire N__3692;
    wire N__3689;
    wire N__3686;
    wire N__3681;
    wire N__3678;
    wire N__3677;
    wire N__3674;
    wire N__3671;
    wire N__3666;
    wire N__3663;
    wire N__3662;
    wire N__3659;
    wire N__3656;
    wire N__3651;
    wire N__3648;
    wire N__3647;
    wire N__3644;
    wire N__3641;
    wire N__3636;
    wire N__3633;
    wire N__3632;
    wire N__3631;
    wire N__3624;
    wire N__3621;
    wire N__3620;
    wire N__3617;
    wire N__3614;
    wire N__3609;
    wire N__3606;
    wire N__3603;
    wire N__3600;
    wire N__3597;
    wire N__3596;
    wire N__3593;
    wire N__3590;
    wire N__3585;
    wire N__3582;
    wire N__3579;
    wire N__3576;
    wire N__3573;
    wire N__3572;
    wire N__3569;
    wire N__3566;
    wire N__3561;
    wire N__3558;
    wire N__3555;
    wire N__3552;
    wire N__3551;
    wire N__3548;
    wire N__3545;
    wire N__3540;
    wire N__3537;
    wire N__3536;
    wire N__3533;
    wire N__3530;
    wire N__3525;
    wire N__3522;
    wire N__3519;
    wire N__3516;
    wire N__3513;
    wire N__3512;
    wire N__3509;
    wire N__3506;
    wire N__3501;
    wire N__3498;
    wire N__3497;
    wire N__3494;
    wire N__3491;
    wire N__3486;
    wire N__3483;
    wire N__3482;
    wire N__3479;
    wire N__3476;
    wire N__3471;
    wire N__3468;
    wire N__3465;
    wire N__3462;
    wire N__3459;
    wire N__3456;
    wire N__3453;
    wire N__3450;
    wire N__3447;
    wire N__3444;
    wire N__3441;
    wire N__3438;
    wire N__3437;
    wire N__3434;
    wire N__3431;
    wire N__3428;
    wire N__3425;
    wire N__3420;
    wire N__3417;
    wire N__3416;
    wire N__3413;
    wire N__3410;
    wire N__3405;
    wire N__3402;
    wire N__3399;
    wire N__3396;
    wire N__3393;
    wire N__3390;
    wire N__3389;
    wire N__3388;
    wire N__3385;
    wire N__3380;
    wire N__3375;
    wire N__3374;
    wire N__3371;
    wire N__3368;
    wire N__3367;
    wire N__3364;
    wire N__3361;
    wire N__3358;
    wire N__3351;
    wire N__3350;
    wire N__3347;
    wire N__3344;
    wire N__3343;
    wire N__3340;
    wire N__3337;
    wire N__3334;
    wire N__3331;
    wire N__3324;
    wire N__3321;
    wire N__3320;
    wire N__3319;
    wire N__3318;
    wire N__3317;
    wire N__3316;
    wire N__3315;
    wire N__3312;
    wire N__3303;
    wire N__3302;
    wire N__3299;
    wire N__3298;
    wire N__3297;
    wire N__3296;
    wire N__3295;
    wire N__3294;
    wire N__3291;
    wire N__3290;
    wire N__3289;
    wire N__3286;
    wire N__3283;
    wire N__3270;
    wire N__3261;
    wire N__3252;
    wire N__3249;
    wire N__3248;
    wire N__3245;
    wire N__3244;
    wire N__3243;
    wire N__3242;
    wire N__3239;
    wire N__3238;
    wire N__3237;
    wire N__3236;
    wire N__3233;
    wire N__3228;
    wire N__3223;
    wire N__3222;
    wire N__3221;
    wire N__3220;
    wire N__3217;
    wire N__3216;
    wire N__3213;
    wire N__3212;
    wire N__3211;
    wire N__3210;
    wire N__3207;
    wire N__3204;
    wire N__3199;
    wire N__3186;
    wire N__3183;
    wire N__3176;
    wire N__3165;
    wire N__3164;
    wire N__3161;
    wire N__3160;
    wire N__3157;
    wire N__3154;
    wire N__3151;
    wire N__3148;
    wire N__3141;
    wire N__3140;
    wire N__3137;
    wire N__3134;
    wire N__3133;
    wire N__3130;
    wire N__3127;
    wire N__3124;
    wire N__3121;
    wire N__3114;
    wire N__3111;
    wire N__3110;
    wire N__3109;
    wire N__3106;
    wire N__3103;
    wire N__3100;
    wire N__3093;
    wire N__3090;
    wire N__3087;
    wire N__3084;
    wire N__3081;
    wire N__3078;
    wire N__3075;
    wire N__3072;
    wire N__3069;
    wire N__3066;
    wire N__3063;
    wire N__3060;
    wire N__3057;
    wire N__3054;
    wire N__3051;
    wire N__3048;
    wire N__3047;
    wire N__3044;
    wire N__3043;
    wire N__3040;
    wire N__3037;
    wire N__3034;
    wire N__3027;
    wire N__3026;
    wire N__3025;
    wire N__3022;
    wire N__3017;
    wire N__3012;
    wire N__3011;
    wire N__3010;
    wire N__3007;
    wire N__3002;
    wire N__2997;
    wire N__2996;
    wire N__2993;
    wire N__2992;
    wire N__2989;
    wire N__2986;
    wire N__2983;
    wire N__2976;
    wire N__2975;
    wire N__2974;
    wire N__2971;
    wire N__2968;
    wire N__2965;
    wire N__2958;
    wire N__2957;
    wire N__2956;
    wire N__2953;
    wire N__2948;
    wire N__2943;
    wire N__2942;
    wire N__2941;
    wire N__2938;
    wire N__2933;
    wire N__2928;
    wire N__2927;
    wire N__2924;
    wire N__2923;
    wire N__2920;
    wire N__2917;
    wire N__2914;
    wire N__2907;
    wire N__2904;
    wire N__2901;
    wire N__2898;
    wire N__2895;
    wire N__2892;
    wire N__2889;
    wire N__2886;
    wire N__2883;
    wire N__2880;
    wire N__2877;
    wire N__2876;
    wire N__2871;
    wire N__2868;
    wire N__2865;
    wire N__2862;
    wire N__2859;
    wire N__2856;
    wire N__2855;
    wire N__2850;
    wire N__2847;
    wire N__2844;
    wire N__2841;
    wire N__2838;
    wire N__2837;
    wire N__2836;
    wire N__2835;
    wire N__2830;
    wire N__2825;
    wire N__2820;
    wire N__2817;
    wire N__2814;
    wire N__2811;
    wire N__2808;
    wire N__2807;
    wire N__2806;
    wire N__2803;
    wire N__2798;
    wire N__2793;
    wire N__2792;
    wire N__2789;
    wire N__2786;
    wire N__2781;
    wire N__2780;
    wire N__2779;
    wire N__2776;
    wire N__2771;
    wire N__2766;
    wire N__2763;
    wire N__2760;
    wire N__2757;
    wire N__2754;
    wire N__2751;
    wire N__2748;
    wire N__2745;
    wire N__2742;
    wire N__2739;
    wire N__2736;
    wire N__2733;
    wire N__2730;
    wire N__2727;
    wire N__2724;
    wire N__2721;
    wire N__2718;
    wire N__2715;
    wire N__2712;
    wire N__2709;
    wire N__2706;
    wire N__2703;
    wire N__2700;
    wire N__2697;
    wire N__2694;
    wire N__2691;
    wire N__2688;
    wire N__2685;
    wire N__2682;
    wire N__2679;
    wire N__2676;
    wire N__2673;
    wire N__2670;
    wire N__2667;
    wire N__2664;
    wire N__2661;
    wire N__2658;
    wire N__2655;
    wire N__2652;
    wire N__2649;
    wire N__2648;
    wire N__2647;
    wire N__2646;
    wire N__2641;
    wire N__2636;
    wire N__2631;
    wire N__2630;
    wire N__2629;
    wire N__2628;
    wire N__2619;
    wire N__2616;
    wire N__2613;
    wire N__2610;
    wire N__2607;
    wire N__2604;
    wire N__2601;
    wire N__2598;
    wire N__2595;
    wire N__2592;
    wire N__2589;
    wire N__2586;
    wire N__2583;
    wire N__2580;
    wire N__2577;
    wire N__2574;
    wire N__2571;
    wire N__2568;
    wire N__2565;
    wire N__2562;
    wire N__2559;
    wire N__2556;
    wire N__2553;
    wire N__2550;
    wire N__2547;
    wire N__2544;
    wire N__2541;
    wire N__2540;
    wire N__2537;
    wire N__2534;
    wire N__2531;
    wire N__2526;
    wire N__2523;
    wire N__2522;
    wire N__2519;
    wire N__2516;
    wire N__2513;
    wire N__2508;
    wire N__2505;
    wire N__2502;
    wire N__2499;
    wire N__2496;
    wire N__2493;
    wire N__2490;
    wire N__2487;
    wire N__2484;
    wire N__2481;
    wire N__2478;
    wire N__2475;
    wire N__2472;
    wire N__2469;
    wire N__2466;
    wire N__2463;
    wire N__2460;
    wire N__2457;
    wire N__2454;
    wire N__2451;
    wire N__2448;
    wire N__2445;
    wire N__2442;
    wire N__2439;
    wire N__2436;
    wire N__2433;
    wire N__2430;
    wire N__2427;
    wire N__2424;
    wire N__2421;
    wire N__2420;
    wire N__2417;
    wire N__2414;
    wire N__2409;
    wire N__2406;
    wire N__2405;
    wire N__2402;
    wire N__2399;
    wire N__2394;
    wire N__2391;
    wire N__2390;
    wire N__2387;
    wire N__2384;
    wire N__2379;
    wire N__2376;
    wire N__2375;
    wire N__2372;
    wire N__2369;
    wire N__2364;
    wire N__2361;
    wire N__2360;
    wire N__2357;
    wire N__2354;
    wire N__2349;
    wire N__2346;
    wire N__2345;
    wire N__2342;
    wire N__2339;
    wire N__2334;
    wire N__2331;
    wire N__2330;
    wire N__2327;
    wire N__2324;
    wire N__2319;
    wire N__2316;
    wire N__2315;
    wire N__2312;
    wire N__2309;
    wire N__2304;
    wire N__2301;
    wire N__2300;
    wire N__2297;
    wire N__2294;
    wire N__2289;
    wire N__2286;
    wire N__2283;
    wire N__2282;
    wire N__2277;
    wire N__2274;
    wire N__2271;
    wire N__2268;
    wire N__2265;
    wire N__2262;
    wire N__2261;
    wire N__2258;
    wire N__2255;
    wire N__2250;
    wire N__2247;
    wire N__2244;
    wire N__2243;
    wire N__2240;
    wire N__2237;
    wire N__2232;
    wire N__2229;
    wire N__2226;
    wire N__2223;
    wire N__2220;
    wire N__2217;
    wire N__2214;
    wire N__2213;
    wire N__2210;
    wire N__2207;
    wire N__2202;
    wire N__2199;
    wire N__2198;
    wire N__2195;
    wire N__2192;
    wire N__2187;
    wire N__2184;
    wire N__2183;
    wire N__2180;
    wire N__2177;
    wire N__2172;
    wire N__2169;
    wire N__2168;
    wire N__2165;
    wire N__2162;
    wire N__2157;
    wire N__2154;
    wire N__2153;
    wire N__2150;
    wire N__2147;
    wire N__2142;
    wire N__2139;
    wire N__2136;
    wire N__2133;
    wire N__2130;
    wire N__2127;
    wire N__2124;
    wire N__2121;
    wire N__2118;
    wire N__2115;
    wire N__2112;
    wire N__2109;
    wire N__2106;
    wire N__2103;
    wire N__2100;
    wire N__2097;
    wire N__2094;
    wire VCCG0;
    wire GNDG0;
    wire bfn_1_7_0_;
    wire \pulse_counter.n728 ;
    wire \pulse_counter.n729 ;
    wire \pulse_counter.n730 ;
    wire \pulse_counter.n731 ;
    wire \pulse_counter.n732 ;
    wire \pulse_counter.n733 ;
    wire \pulse_counter.n734 ;
    wire \pulse_counter.n735 ;
    wire bfn_1_8_0_;
    wire \pulse_counter.n736 ;
    wire \pulse_counter.n737 ;
    wire \pulse_counter.n738 ;
    wire \pulse_counter.n739 ;
    wire \pulse_counter.n740 ;
    wire \pulse_counter.n741 ;
    wire \pulse_counter.n742 ;
    wire divide_enable_c;
    wire n176;
    wire output_state;
    wire constant_v_c;
    wire \pulse_counter.internal_count_0 ;
    wire bfn_2_7_0_;
    wire \pulse_counter.internal_count_1 ;
    wire \pulse_counter.n712 ;
    wire \pulse_counter.internal_count_2 ;
    wire \pulse_counter.n713 ;
    wire \pulse_counter.internal_count_3 ;
    wire \pulse_counter.n714 ;
    wire \pulse_counter.internal_count_4 ;
    wire \pulse_counter.n715 ;
    wire \pulse_counter.internal_count_5 ;
    wire \pulse_counter.n716 ;
    wire \pulse_counter.internal_count_6 ;
    wire \pulse_counter.n717 ;
    wire \pulse_counter.internal_count_7 ;
    wire \pulse_counter.n718 ;
    wire \pulse_counter.n719 ;
    wire \pulse_counter.internal_count_8 ;
    wire bfn_2_8_0_;
    wire \pulse_counter.internal_count_9 ;
    wire \pulse_counter.n720 ;
    wire \pulse_counter.internal_count_10 ;
    wire \pulse_counter.n721 ;
    wire \pulse_counter.internal_count_11 ;
    wire \pulse_counter.n722 ;
    wire \pulse_counter.internal_count_12 ;
    wire \pulse_counter.n723 ;
    wire \pulse_counter.internal_count_13 ;
    wire \pulse_counter.n724 ;
    wire \pulse_counter.internal_count_14 ;
    wire \pulse_counter.n725 ;
    wire \pulse_counter.internal_count_15 ;
    wire \pulse_counter.n726 ;
    wire \pulse_counter.n727 ;
    wire \pulse_counter.n13 ;
    wire bfn_2_9_0_;
    wire n4_adj_116;
    wire n5_adj_120;
    wire n1_adj_117;
    wire n9;
    wire n795_cascade_;
    wire n6_adj_119;
    wire n12;
    wire n16;
    wire n817_cascade_;
    wire n787;
    wire n825_cascade_;
    wire sr_divider_data_11;
    wire sr_divider_data_13;
    wire count_done;
    wire laser_pulse_c;
    wire sr_divider_data_2;
    wire sr_divider_data_14;
    wire sr_divider_data_15;
    wire sr_divider_data_0;
    wire sr_divider_data_3;
    wire sr_divider_data_12;
    wire sr_divider_data_1;
    wire sr_divider_data_10;
    wire sr_divider_data_6;
    wire sr_divider_data_9;
    wire sr_divider_data_4;
    wire sr_divider_data_5;
    wire sr_divider_data_8;
    wire sr_divider_data_7;
    wire n8;
    wire n3_adj_118;
    wire n15;
    wire n7;
    wire n10;
    wire n14;
    wire n2_adj_99;
    wire n11;
    wire n823_cascade_;
    wire n781;
    wire n827;
    wire sr_sel_row_c;
    wire n169_cascade_;
    wire sr_sel_div_c;
    wire sr_reset_c;
    wire n330_cascade_;
    wire shifted_data_14;
    wire shifted_data_15;
    wire shifted_data_11;
    wire shifted_data_12;
    wire shifted_data_13;
    wire shifted_data_8;
    wire shifted_data_9;
    wire shifted_data_10;
    wire shifted_data_5;
    wire shifted_data_6;
    wire shifted_data_7;
    wire bfn_5_7_0_;
    wire \row_counter.n743 ;
    wire \row_counter.n744 ;
    wire \row_counter.n745 ;
    wire \row_counter.n746 ;
    wire \row_counter.n747 ;
    wire \row_counter.n748 ;
    wire \row_counter.n749 ;
    wire \row_counter.n750 ;
    wire bfn_5_8_0_;
    wire \row_counter.n751 ;
    wire \row_counter.n752 ;
    wire \row_counter.n753 ;
    wire \row_counter.n754 ;
    wire \row_counter.n755 ;
    wire \row_counter.n756 ;
    wire \row_counter.n757 ;
    wire en_rowpack_c;
    wire n189;
    wire sr_data_c;
    wire shifted_data_0;
    wire shifted_data_1;
    wire shifted_data_2;
    wire n330;
    wire n169;
    wire shifted_data_3;
    wire shifted_data_4;
    wire shifted_data_0_adj_115;
    wire shifted_data_1_adj_114;
    wire \row_counter.internal_count_0 ;
    wire sr_row_data_0;
    wire bfn_6_7_0_;
    wire \row_counter.internal_count_1 ;
    wire sr_row_data_1;
    wire \row_counter.n696 ;
    wire \row_counter.internal_count_2 ;
    wire \row_counter.n697 ;
    wire \row_counter.internal_count_3 ;
    wire \row_counter.n698 ;
    wire \row_counter.internal_count_4 ;
    wire sr_row_data_4;
    wire \row_counter.n699 ;
    wire \row_counter.internal_count_5 ;
    wire \row_counter.n700 ;
    wire \row_counter.internal_count_6 ;
    wire \row_counter.n701 ;
    wire \row_counter.internal_count_7 ;
    wire sr_row_data_7;
    wire \row_counter.n702 ;
    wire \row_counter.n703 ;
    wire \row_counter.internal_count_8 ;
    wire bfn_6_8_0_;
    wire \row_counter.internal_count_9 ;
    wire \row_counter.n704 ;
    wire \row_counter.internal_count_10 ;
    wire \row_counter.n705 ;
    wire \row_counter.internal_count_11 ;
    wire \row_counter.n706 ;
    wire \row_counter.internal_count_12 ;
    wire \row_counter.n707 ;
    wire \row_counter.internal_count_13 ;
    wire \row_counter.n708 ;
    wire \row_counter.internal_count_14 ;
    wire \row_counter.n709 ;
    wire \row_counter.internal_count_15 ;
    wire \row_counter.n710 ;
    wire \row_counter.n711 ;
    wire \row_counter.n13 ;
    wire CONSTANT_ONE_NET;
    wire bfn_6_9_0_;
    wire sr_row_data_8;
    wire sr_row_data_6;
    wire sr_row_data_9;
    wire n4;
    wire n5;
    wire n1;
    wire n9_adj_123;
    wire n811_cascade_;
    wire n6;
    wire n12_adj_126;
    wire n16_adj_129;
    wire n831_cascade_;
    wire n775;
    wire reset_signal;
    wire n835_cascade_;
    wire row_complete;
    wire divided_pulse_c;
    wire sr_row_data_14;
    wire sr_row_data_11;
    wire sr_row_data_15;
    wire sr_row_data_13;
    wire shifted_data_15_adj_100;
    wire shifted_data_14_adj_101;
    wire sr_row_data_10;
    wire shifted_data_2_adj_113;
    wire sr_row_data_2;
    wire n8_adj_122;
    wire n3;
    wire shifted_data_4_adj_111;
    wire n15_adj_128;
    wire n7_adj_121;
    wire n10_adj_124;
    wire n14_adj_127;
    wire n2;
    wire n11_adj_125;
    wire n793_cascade_;
    wire n803;
    wire n829;
    wire shifted_data_6_adj_109;
    wire shifted_data_7_adj_108;
    wire shifted_data_8_adj_107;
    wire sr_row_data_12;
    wire shifted_data_13_adj_102;
    wire shifted_data_11_adj_104;
    wire shifted_data_12_adj_103;
    wire n345;
    wire n171;
    wire shifted_data_9_adj_106;
    wire shifted_data_10_adj_105;
    wire sr_clk_c;
    wire shifted_data_5_adj_110;
    wire sr_row_data_5;
    wire en_internals_c;
    wire shifted_data_3_adj_112;
    wire sr_row_data_3;
    wire _gnd_net_;

    PRE_IO_GBUF sr_clk_pad_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__5168),
            .GLOBALBUFFEROUTPUT(sr_clk_c));
    defparam sr_clk_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam sr_clk_pad_iopad.PULLUP=1'b0;
    IO_PAD sr_clk_pad_iopad (
            .OE(N__5170),
            .DIN(N__5169),
            .DOUT(N__5168),
            .PACKAGEPIN(sr_clk));
    defparam sr_clk_pad_preio.PIN_TYPE=6'b000001;
    defparam sr_clk_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO sr_clk_pad_preio (
            .PADOEN(N__5170),
            .PADOUT(N__5169),
            .PADIN(N__5168),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF laser_pulse_pad_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__5158),
            .GLOBALBUFFEROUTPUT(laser_pulse_c));
    defparam laser_pulse_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam laser_pulse_pad_iopad.PULLUP=1'b0;
    IO_PAD laser_pulse_pad_iopad (
            .OE(N__5160),
            .DIN(N__5159),
            .DOUT(N__5158),
            .PACKAGEPIN(laser_pulse));
    defparam laser_pulse_pad_preio.PIN_TYPE=6'b000001;
    defparam laser_pulse_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO laser_pulse_pad_preio (
            .PADOEN(N__5160),
            .PADOUT(N__5159),
            .PADIN(N__5158),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam en_internals_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam en_internals_pad_iopad.PULLUP=1'b0;
    IO_PAD en_internals_pad_iopad (
            .OE(N__5149),
            .DIN(N__5148),
            .DOUT(N__5147),
            .PACKAGEPIN(en_internals));
    defparam en_internals_pad_preio.PIN_TYPE=6'b000001;
    defparam en_internals_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO en_internals_pad_preio (
            .PADOEN(N__5149),
            .PADOUT(N__5148),
            .PADIN(N__5147),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(en_internals_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam sr_reset_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam sr_reset_pad_iopad.PULLUP=1'b0;
    IO_PAD sr_reset_pad_iopad (
            .OE(N__5140),
            .DIN(N__5139),
            .DOUT(N__5138),
            .PACKAGEPIN(sr_reset));
    defparam sr_reset_pad_preio.PIN_TYPE=6'b000001;
    defparam sr_reset_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO sr_reset_pad_preio (
            .PADOEN(N__5140),
            .PADOUT(N__5139),
            .PADIN(N__5138),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(sr_reset_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam sr_data_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam sr_data_pad_iopad.PULLUP=1'b0;
    IO_PAD sr_data_pad_iopad (
            .OE(N__5131),
            .DIN(N__5130),
            .DOUT(N__5129),
            .PACKAGEPIN(sr_data));
    defparam sr_data_pad_preio.PIN_TYPE=6'b000001;
    defparam sr_data_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO sr_data_pad_preio (
            .PADOEN(N__5131),
            .PADOUT(N__5130),
            .PADIN(N__5129),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(sr_data_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam divide_enable_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam divide_enable_pad_iopad.PULLUP=1'b0;
    IO_PAD divide_enable_pad_iopad (
            .OE(N__5122),
            .DIN(N__5121),
            .DOUT(N__5120),
            .PACKAGEPIN(divide_enable));
    defparam divide_enable_pad_preio.PIN_TYPE=6'b000001;
    defparam divide_enable_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO divide_enable_pad_preio (
            .PADOEN(N__5122),
            .PADOUT(N__5121),
            .PADIN(N__5120),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(divide_enable_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam sr_sel_div_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam sr_sel_div_pad_iopad.PULLUP=1'b0;
    IO_PAD sr_sel_div_pad_iopad (
            .OE(N__5113),
            .DIN(N__5112),
            .DOUT(N__5111),
            .PACKAGEPIN(sr_sel_div));
    defparam sr_sel_div_pad_preio.PIN_TYPE=6'b000001;
    defparam sr_sel_div_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO sr_sel_div_pad_preio (
            .PADOEN(N__5113),
            .PADOUT(N__5112),
            .PADIN(N__5111),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(sr_sel_div_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam constant_v_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam constant_v_pad_iopad.PULLUP=1'b0;
    IO_PAD constant_v_pad_iopad (
            .OE(N__5104),
            .DIN(N__5103),
            .DOUT(N__5102),
            .PACKAGEPIN(constant_v));
    defparam constant_v_pad_preio.PIN_TYPE=6'b000001;
    defparam constant_v_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO constant_v_pad_preio (
            .PADOEN(N__5104),
            .PADOUT(N__5103),
            .PADIN(N__5102),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(constant_v_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam divided_pulse_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam divided_pulse_pad_iopad.PULLUP=1'b0;
    IO_PAD divided_pulse_pad_iopad (
            .OE(N__5095),
            .DIN(N__5094),
            .DOUT(N__5093),
            .PACKAGEPIN(divided_pulse));
    defparam divided_pulse_pad_preio.PIN_TYPE=6'b011001;
    defparam divided_pulse_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO divided_pulse_pad_preio (
            .PADOEN(N__5095),
            .PADOUT(N__5094),
            .PADIN(N__5093),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3789),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam en_rowpack_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam en_rowpack_pad_iopad.PULLUP=1'b0;
    IO_PAD en_rowpack_pad_iopad (
            .OE(N__5086),
            .DIN(N__5085),
            .DOUT(N__5084),
            .PACKAGEPIN(en_rowpack));
    defparam en_rowpack_pad_preio.PIN_TYPE=6'b000001;
    defparam en_rowpack_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO en_rowpack_pad_preio (
            .PADOEN(N__5086),
            .PADOUT(N__5085),
            .PADIN(N__5084),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(en_rowpack_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam sr_sel_row_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam sr_sel_row_pad_iopad.PULLUP=1'b0;
    IO_PAD sr_sel_row_pad_iopad (
            .OE(N__5077),
            .DIN(N__5076),
            .DOUT(N__5075),
            .PACKAGEPIN(sr_sel_row));
    defparam sr_sel_row_pad_preio.PIN_TYPE=6'b000001;
    defparam sr_sel_row_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO sr_sel_row_pad_preio (
            .PADOEN(N__5077),
            .PADOUT(N__5076),
            .PADIN(N__5075),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(sr_sel_row_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam row_completed_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam row_completed_pad_iopad.PULLUP=1'b0;
    IO_PAD row_completed_pad_iopad (
            .OE(N__5068),
            .DIN(N__5067),
            .DOUT(N__5066),
            .PACKAGEPIN(row_completed));
    defparam row_completed_pad_preio.PIN_TYPE=6'b011001;
    defparam row_completed_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO row_completed_pad_preio (
            .PADOEN(N__5068),
            .PADOUT(N__5067),
            .PADIN(N__5066),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1164 (
            .O(N__5049),
            .I(N__5044));
    InMux I__1163 (
            .O(N__5048),
            .I(N__5039));
    InMux I__1162 (
            .O(N__5047),
            .I(N__5039));
    LocalMux I__1161 (
            .O(N__5044),
            .I(shifted_data_8_adj_107));
    LocalMux I__1160 (
            .O(N__5039),
            .I(shifted_data_8_adj_107));
    InMux I__1159 (
            .O(N__5034),
            .I(N__5031));
    LocalMux I__1158 (
            .O(N__5031),
            .I(N__5028));
    Odrv4 I__1157 (
            .O(N__5028),
            .I(sr_row_data_12));
    CascadeMux I__1156 (
            .O(N__5025),
            .I(N__5020));
    InMux I__1155 (
            .O(N__5024),
            .I(N__5015));
    InMux I__1154 (
            .O(N__5023),
            .I(N__5015));
    InMux I__1153 (
            .O(N__5020),
            .I(N__5012));
    LocalMux I__1152 (
            .O(N__5015),
            .I(shifted_data_13_adj_102));
    LocalMux I__1151 (
            .O(N__5012),
            .I(shifted_data_13_adj_102));
    CascadeMux I__1150 (
            .O(N__5007),
            .I(N__5004));
    InMux I__1149 (
            .O(N__5004),
            .I(N__4999));
    InMux I__1148 (
            .O(N__5003),
            .I(N__4994));
    InMux I__1147 (
            .O(N__5002),
            .I(N__4994));
    LocalMux I__1146 (
            .O(N__4999),
            .I(shifted_data_11_adj_104));
    LocalMux I__1145 (
            .O(N__4994),
            .I(shifted_data_11_adj_104));
    InMux I__1144 (
            .O(N__4989),
            .I(N__4980));
    InMux I__1143 (
            .O(N__4988),
            .I(N__4980));
    InMux I__1142 (
            .O(N__4987),
            .I(N__4980));
    LocalMux I__1141 (
            .O(N__4980),
            .I(shifted_data_12_adj_103));
    CascadeMux I__1140 (
            .O(N__4977),
            .I(N__4972));
    InMux I__1139 (
            .O(N__4976),
            .I(N__4958));
    InMux I__1138 (
            .O(N__4975),
            .I(N__4951));
    InMux I__1137 (
            .O(N__4972),
            .I(N__4951));
    InMux I__1136 (
            .O(N__4971),
            .I(N__4951));
    InMux I__1135 (
            .O(N__4970),
            .I(N__4948));
    InMux I__1134 (
            .O(N__4969),
            .I(N__4941));
    InMux I__1133 (
            .O(N__4968),
            .I(N__4941));
    InMux I__1132 (
            .O(N__4967),
            .I(N__4941));
    InMux I__1131 (
            .O(N__4966),
            .I(N__4936));
    InMux I__1130 (
            .O(N__4965),
            .I(N__4936));
    InMux I__1129 (
            .O(N__4964),
            .I(N__4933));
    InMux I__1128 (
            .O(N__4963),
            .I(N__4926));
    InMux I__1127 (
            .O(N__4962),
            .I(N__4926));
    InMux I__1126 (
            .O(N__4961),
            .I(N__4926));
    LocalMux I__1125 (
            .O(N__4958),
            .I(N__4917));
    LocalMux I__1124 (
            .O(N__4951),
            .I(N__4917));
    LocalMux I__1123 (
            .O(N__4948),
            .I(N__4917));
    LocalMux I__1122 (
            .O(N__4941),
            .I(N__4914));
    LocalMux I__1121 (
            .O(N__4936),
            .I(N__4909));
    LocalMux I__1120 (
            .O(N__4933),
            .I(N__4909));
    LocalMux I__1119 (
            .O(N__4926),
            .I(N__4906));
    InMux I__1118 (
            .O(N__4925),
            .I(N__4901));
    InMux I__1117 (
            .O(N__4924),
            .I(N__4901));
    Span4Mux_v I__1116 (
            .O(N__4917),
            .I(N__4896));
    Span4Mux_v I__1115 (
            .O(N__4914),
            .I(N__4896));
    Span4Mux_v I__1114 (
            .O(N__4909),
            .I(N__4891));
    Span4Mux_v I__1113 (
            .O(N__4906),
            .I(N__4891));
    LocalMux I__1112 (
            .O(N__4901),
            .I(N__4888));
    Odrv4 I__1111 (
            .O(N__4896),
            .I(n345));
    Odrv4 I__1110 (
            .O(N__4891),
            .I(n345));
    Odrv12 I__1109 (
            .O(N__4888),
            .I(n345));
    CascadeMux I__1108 (
            .O(N__4881),
            .I(N__4873));
    CascadeMux I__1107 (
            .O(N__4880),
            .I(N__4868));
    CascadeMux I__1106 (
            .O(N__4879),
            .I(N__4865));
    CascadeMux I__1105 (
            .O(N__4878),
            .I(N__4859));
    CascadeMux I__1104 (
            .O(N__4877),
            .I(N__4856));
    CascadeMux I__1103 (
            .O(N__4876),
            .I(N__4853));
    InMux I__1102 (
            .O(N__4873),
            .I(N__4846));
    InMux I__1101 (
            .O(N__4872),
            .I(N__4846));
    InMux I__1100 (
            .O(N__4871),
            .I(N__4846));
    InMux I__1099 (
            .O(N__4868),
            .I(N__4841));
    InMux I__1098 (
            .O(N__4865),
            .I(N__4841));
    CascadeMux I__1097 (
            .O(N__4864),
            .I(N__4836));
    CascadeMux I__1096 (
            .O(N__4863),
            .I(N__4832));
    CascadeMux I__1095 (
            .O(N__4862),
            .I(N__4829));
    InMux I__1094 (
            .O(N__4859),
            .I(N__4825));
    InMux I__1093 (
            .O(N__4856),
            .I(N__4822));
    InMux I__1092 (
            .O(N__4853),
            .I(N__4819));
    LocalMux I__1091 (
            .O(N__4846),
            .I(N__4814));
    LocalMux I__1090 (
            .O(N__4841),
            .I(N__4814));
    InMux I__1089 (
            .O(N__4840),
            .I(N__4809));
    InMux I__1088 (
            .O(N__4839),
            .I(N__4809));
    InMux I__1087 (
            .O(N__4836),
            .I(N__4806));
    InMux I__1086 (
            .O(N__4835),
            .I(N__4799));
    InMux I__1085 (
            .O(N__4832),
            .I(N__4799));
    InMux I__1084 (
            .O(N__4829),
            .I(N__4799));
    CascadeMux I__1083 (
            .O(N__4828),
            .I(N__4795));
    LocalMux I__1082 (
            .O(N__4825),
            .I(N__4792));
    LocalMux I__1081 (
            .O(N__4822),
            .I(N__4787));
    LocalMux I__1080 (
            .O(N__4819),
            .I(N__4787));
    Span4Mux_v I__1079 (
            .O(N__4814),
            .I(N__4778));
    LocalMux I__1078 (
            .O(N__4809),
            .I(N__4778));
    LocalMux I__1077 (
            .O(N__4806),
            .I(N__4778));
    LocalMux I__1076 (
            .O(N__4799),
            .I(N__4778));
    InMux I__1075 (
            .O(N__4798),
            .I(N__4773));
    InMux I__1074 (
            .O(N__4795),
            .I(N__4773));
    Span4Mux_v I__1073 (
            .O(N__4792),
            .I(N__4770));
    Span4Mux_v I__1072 (
            .O(N__4787),
            .I(N__4765));
    Span4Mux_v I__1071 (
            .O(N__4778),
            .I(N__4765));
    LocalMux I__1070 (
            .O(N__4773),
            .I(N__4762));
    Odrv4 I__1069 (
            .O(N__4770),
            .I(n171));
    Odrv4 I__1068 (
            .O(N__4765),
            .I(n171));
    Odrv12 I__1067 (
            .O(N__4762),
            .I(n171));
    CascadeMux I__1066 (
            .O(N__4755),
            .I(N__4750));
    InMux I__1065 (
            .O(N__4754),
            .I(N__4747));
    InMux I__1064 (
            .O(N__4753),
            .I(N__4744));
    InMux I__1063 (
            .O(N__4750),
            .I(N__4741));
    LocalMux I__1062 (
            .O(N__4747),
            .I(shifted_data_9_adj_106));
    LocalMux I__1061 (
            .O(N__4744),
            .I(shifted_data_9_adj_106));
    LocalMux I__1060 (
            .O(N__4741),
            .I(shifted_data_9_adj_106));
    InMux I__1059 (
            .O(N__4734),
            .I(N__4727));
    InMux I__1058 (
            .O(N__4733),
            .I(N__4727));
    InMux I__1057 (
            .O(N__4732),
            .I(N__4724));
    LocalMux I__1056 (
            .O(N__4727),
            .I(shifted_data_10_adj_105));
    LocalMux I__1055 (
            .O(N__4724),
            .I(shifted_data_10_adj_105));
    ClkMux I__1054 (
            .O(N__4719),
            .I(N__4683));
    ClkMux I__1053 (
            .O(N__4718),
            .I(N__4683));
    ClkMux I__1052 (
            .O(N__4717),
            .I(N__4683));
    ClkMux I__1051 (
            .O(N__4716),
            .I(N__4683));
    ClkMux I__1050 (
            .O(N__4715),
            .I(N__4683));
    ClkMux I__1049 (
            .O(N__4714),
            .I(N__4683));
    ClkMux I__1048 (
            .O(N__4713),
            .I(N__4683));
    ClkMux I__1047 (
            .O(N__4712),
            .I(N__4683));
    ClkMux I__1046 (
            .O(N__4711),
            .I(N__4683));
    ClkMux I__1045 (
            .O(N__4710),
            .I(N__4683));
    ClkMux I__1044 (
            .O(N__4709),
            .I(N__4683));
    ClkMux I__1043 (
            .O(N__4708),
            .I(N__4683));
    GlobalMux I__1042 (
            .O(N__4683),
            .I(N__4680));
    gio2CtrlBuf I__1041 (
            .O(N__4680),
            .I(sr_clk_c));
    InMux I__1040 (
            .O(N__4677),
            .I(N__4672));
    InMux I__1039 (
            .O(N__4676),
            .I(N__4667));
    InMux I__1038 (
            .O(N__4675),
            .I(N__4667));
    LocalMux I__1037 (
            .O(N__4672),
            .I(shifted_data_5_adj_110));
    LocalMux I__1036 (
            .O(N__4667),
            .I(shifted_data_5_adj_110));
    CascadeMux I__1035 (
            .O(N__4662),
            .I(N__4659));
    InMux I__1034 (
            .O(N__4659),
            .I(N__4656));
    LocalMux I__1033 (
            .O(N__4656),
            .I(N__4653));
    Odrv4 I__1032 (
            .O(N__4653),
            .I(sr_row_data_5));
    InMux I__1031 (
            .O(N__4650),
            .I(N__4642));
    InMux I__1030 (
            .O(N__4649),
            .I(N__4639));
    InMux I__1029 (
            .O(N__4648),
            .I(N__4632));
    InMux I__1028 (
            .O(N__4647),
            .I(N__4632));
    InMux I__1027 (
            .O(N__4646),
            .I(N__4632));
    InMux I__1026 (
            .O(N__4645),
            .I(N__4624));
    LocalMux I__1025 (
            .O(N__4642),
            .I(N__4612));
    LocalMux I__1024 (
            .O(N__4639),
            .I(N__4612));
    LocalMux I__1023 (
            .O(N__4632),
            .I(N__4612));
    InMux I__1022 (
            .O(N__4631),
            .I(N__4601));
    InMux I__1021 (
            .O(N__4630),
            .I(N__4601));
    InMux I__1020 (
            .O(N__4629),
            .I(N__4601));
    InMux I__1019 (
            .O(N__4628),
            .I(N__4601));
    InMux I__1018 (
            .O(N__4627),
            .I(N__4601));
    LocalMux I__1017 (
            .O(N__4624),
            .I(N__4598));
    InMux I__1016 (
            .O(N__4623),
            .I(N__4593));
    InMux I__1015 (
            .O(N__4622),
            .I(N__4593));
    InMux I__1014 (
            .O(N__4621),
            .I(N__4578));
    InMux I__1013 (
            .O(N__4620),
            .I(N__4578));
    InMux I__1012 (
            .O(N__4619),
            .I(N__4578));
    Span4Mux_v I__1011 (
            .O(N__4612),
            .I(N__4573));
    LocalMux I__1010 (
            .O(N__4601),
            .I(N__4573));
    Span4Mux_h I__1009 (
            .O(N__4598),
            .I(N__4568));
    LocalMux I__1008 (
            .O(N__4593),
            .I(N__4568));
    InMux I__1007 (
            .O(N__4592),
            .I(N__4551));
    InMux I__1006 (
            .O(N__4591),
            .I(N__4551));
    InMux I__1005 (
            .O(N__4590),
            .I(N__4551));
    InMux I__1004 (
            .O(N__4589),
            .I(N__4551));
    InMux I__1003 (
            .O(N__4588),
            .I(N__4551));
    InMux I__1002 (
            .O(N__4587),
            .I(N__4551));
    InMux I__1001 (
            .O(N__4586),
            .I(N__4551));
    InMux I__1000 (
            .O(N__4585),
            .I(N__4551));
    LocalMux I__999 (
            .O(N__4578),
            .I(N__4540));
    Span4Mux_h I__998 (
            .O(N__4573),
            .I(N__4533));
    Span4Mux_v I__997 (
            .O(N__4568),
            .I(N__4533));
    LocalMux I__996 (
            .O(N__4551),
            .I(N__4533));
    InMux I__995 (
            .O(N__4550),
            .I(N__4520));
    InMux I__994 (
            .O(N__4549),
            .I(N__4520));
    InMux I__993 (
            .O(N__4548),
            .I(N__4520));
    InMux I__992 (
            .O(N__4547),
            .I(N__4520));
    InMux I__991 (
            .O(N__4546),
            .I(N__4520));
    InMux I__990 (
            .O(N__4545),
            .I(N__4520));
    InMux I__989 (
            .O(N__4544),
            .I(N__4515));
    InMux I__988 (
            .O(N__4543),
            .I(N__4515));
    Span4Mux_v I__987 (
            .O(N__4540),
            .I(N__4512));
    Span4Mux_h I__986 (
            .O(N__4533),
            .I(N__4507));
    LocalMux I__985 (
            .O(N__4520),
            .I(N__4507));
    LocalMux I__984 (
            .O(N__4515),
            .I(N__4504));
    Span4Mux_v I__983 (
            .O(N__4512),
            .I(N__4501));
    Span4Mux_v I__982 (
            .O(N__4507),
            .I(N__4498));
    Span12Mux_v I__981 (
            .O(N__4504),
            .I(N__4491));
    Sp12to4 I__980 (
            .O(N__4501),
            .I(N__4491));
    Sp12to4 I__979 (
            .O(N__4498),
            .I(N__4491));
    Odrv12 I__978 (
            .O(N__4491),
            .I(en_internals_c));
    CascadeMux I__977 (
            .O(N__4488),
            .I(N__4485));
    InMux I__976 (
            .O(N__4485),
            .I(N__4481));
    InMux I__975 (
            .O(N__4484),
            .I(N__4477));
    LocalMux I__974 (
            .O(N__4481),
            .I(N__4474));
    InMux I__973 (
            .O(N__4480),
            .I(N__4471));
    LocalMux I__972 (
            .O(N__4477),
            .I(shifted_data_3_adj_112));
    Odrv4 I__971 (
            .O(N__4474),
            .I(shifted_data_3_adj_112));
    LocalMux I__970 (
            .O(N__4471),
            .I(shifted_data_3_adj_112));
    CascadeMux I__969 (
            .O(N__4464),
            .I(N__4461));
    InMux I__968 (
            .O(N__4461),
            .I(N__4458));
    LocalMux I__967 (
            .O(N__4458),
            .I(N__4455));
    Odrv4 I__966 (
            .O(N__4455),
            .I(sr_row_data_3));
    InMux I__965 (
            .O(N__4452),
            .I(N__4447));
    InMux I__964 (
            .O(N__4451),
            .I(N__4444));
    InMux I__963 (
            .O(N__4450),
            .I(N__4441));
    LocalMux I__962 (
            .O(N__4447),
            .I(shifted_data_2_adj_113));
    LocalMux I__961 (
            .O(N__4444),
            .I(shifted_data_2_adj_113));
    LocalMux I__960 (
            .O(N__4441),
            .I(shifted_data_2_adj_113));
    InMux I__959 (
            .O(N__4434),
            .I(N__4431));
    LocalMux I__958 (
            .O(N__4431),
            .I(sr_row_data_2));
    InMux I__957 (
            .O(N__4428),
            .I(N__4425));
    LocalMux I__956 (
            .O(N__4425),
            .I(n8_adj_122));
    InMux I__955 (
            .O(N__4422),
            .I(N__4419));
    LocalMux I__954 (
            .O(N__4419),
            .I(n3));
    InMux I__953 (
            .O(N__4416),
            .I(N__4413));
    LocalMux I__952 (
            .O(N__4413),
            .I(N__4410));
    Span4Mux_v I__951 (
            .O(N__4410),
            .I(N__4405));
    InMux I__950 (
            .O(N__4409),
            .I(N__4400));
    InMux I__949 (
            .O(N__4408),
            .I(N__4400));
    Odrv4 I__948 (
            .O(N__4405),
            .I(shifted_data_4_adj_111));
    LocalMux I__947 (
            .O(N__4400),
            .I(shifted_data_4_adj_111));
    InMux I__946 (
            .O(N__4395),
            .I(N__4392));
    LocalMux I__945 (
            .O(N__4392),
            .I(n15_adj_128));
    InMux I__944 (
            .O(N__4389),
            .I(N__4386));
    LocalMux I__943 (
            .O(N__4386),
            .I(n7_adj_121));
    CascadeMux I__942 (
            .O(N__4383),
            .I(N__4380));
    InMux I__941 (
            .O(N__4380),
            .I(N__4377));
    LocalMux I__940 (
            .O(N__4377),
            .I(n10_adj_124));
    InMux I__939 (
            .O(N__4374),
            .I(N__4371));
    LocalMux I__938 (
            .O(N__4371),
            .I(n14_adj_127));
    InMux I__937 (
            .O(N__4368),
            .I(N__4365));
    LocalMux I__936 (
            .O(N__4365),
            .I(n2));
    InMux I__935 (
            .O(N__4362),
            .I(N__4359));
    LocalMux I__934 (
            .O(N__4359),
            .I(n11_adj_125));
    CascadeMux I__933 (
            .O(N__4356),
            .I(n793_cascade_));
    InMux I__932 (
            .O(N__4353),
            .I(N__4350));
    LocalMux I__931 (
            .O(N__4350),
            .I(n803));
    InMux I__930 (
            .O(N__4347),
            .I(N__4344));
    LocalMux I__929 (
            .O(N__4344),
            .I(n829));
    InMux I__928 (
            .O(N__4341),
            .I(N__4338));
    LocalMux I__927 (
            .O(N__4338),
            .I(N__4333));
    InMux I__926 (
            .O(N__4337),
            .I(N__4330));
    InMux I__925 (
            .O(N__4336),
            .I(N__4327));
    Odrv4 I__924 (
            .O(N__4333),
            .I(shifted_data_6_adj_109));
    LocalMux I__923 (
            .O(N__4330),
            .I(shifted_data_6_adj_109));
    LocalMux I__922 (
            .O(N__4327),
            .I(shifted_data_6_adj_109));
    InMux I__921 (
            .O(N__4320),
            .I(N__4317));
    LocalMux I__920 (
            .O(N__4317),
            .I(N__4314));
    Span4Mux_v I__919 (
            .O(N__4314),
            .I(N__4309));
    InMux I__918 (
            .O(N__4313),
            .I(N__4306));
    InMux I__917 (
            .O(N__4312),
            .I(N__4303));
    Odrv4 I__916 (
            .O(N__4309),
            .I(shifted_data_7_adj_108));
    LocalMux I__915 (
            .O(N__4306),
            .I(shifted_data_7_adj_108));
    LocalMux I__914 (
            .O(N__4303),
            .I(shifted_data_7_adj_108));
    InMux I__913 (
            .O(N__4296),
            .I(N__4293));
    LocalMux I__912 (
            .O(N__4293),
            .I(N__4290));
    Odrv4 I__911 (
            .O(N__4290),
            .I(sr_row_data_14));
    InMux I__910 (
            .O(N__4287),
            .I(N__4284));
    LocalMux I__909 (
            .O(N__4284),
            .I(N__4281));
    Odrv4 I__908 (
            .O(N__4281),
            .I(sr_row_data_11));
    InMux I__907 (
            .O(N__4278),
            .I(N__4275));
    LocalMux I__906 (
            .O(N__4275),
            .I(N__4272));
    Odrv4 I__905 (
            .O(N__4272),
            .I(sr_row_data_15));
    InMux I__904 (
            .O(N__4269),
            .I(N__4266));
    LocalMux I__903 (
            .O(N__4266),
            .I(N__4263));
    Odrv4 I__902 (
            .O(N__4263),
            .I(sr_row_data_13));
    CascadeMux I__901 (
            .O(N__4260),
            .I(N__4256));
    InMux I__900 (
            .O(N__4259),
            .I(N__4251));
    InMux I__899 (
            .O(N__4256),
            .I(N__4251));
    LocalMux I__898 (
            .O(N__4251),
            .I(shifted_data_15_adj_100));
    InMux I__897 (
            .O(N__4248),
            .I(N__4239));
    InMux I__896 (
            .O(N__4247),
            .I(N__4239));
    InMux I__895 (
            .O(N__4246),
            .I(N__4239));
    LocalMux I__894 (
            .O(N__4239),
            .I(shifted_data_14_adj_101));
    InMux I__893 (
            .O(N__4236),
            .I(N__4233));
    LocalMux I__892 (
            .O(N__4233),
            .I(N__4230));
    Odrv4 I__891 (
            .O(N__4230),
            .I(sr_row_data_10));
    InMux I__890 (
            .O(N__4227),
            .I(N__4224));
    LocalMux I__889 (
            .O(N__4224),
            .I(\row_counter.n13 ));
    CascadeMux I__888 (
            .O(N__4221),
            .I(N__4209));
    CascadeMux I__887 (
            .O(N__4220),
            .I(N__4206));
    CascadeMux I__886 (
            .O(N__4219),
            .I(N__4202));
    CascadeMux I__885 (
            .O(N__4218),
            .I(N__4198));
    CascadeMux I__884 (
            .O(N__4217),
            .I(N__4194));
    CascadeMux I__883 (
            .O(N__4216),
            .I(N__4191));
    CascadeMux I__882 (
            .O(N__4215),
            .I(N__4186));
    CascadeMux I__881 (
            .O(N__4214),
            .I(N__4183));
    CascadeMux I__880 (
            .O(N__4213),
            .I(N__4180));
    CascadeMux I__879 (
            .O(N__4212),
            .I(N__4177));
    InMux I__878 (
            .O(N__4209),
            .I(N__4164));
    InMux I__877 (
            .O(N__4206),
            .I(N__4164));
    InMux I__876 (
            .O(N__4205),
            .I(N__4164));
    InMux I__875 (
            .O(N__4202),
            .I(N__4164));
    InMux I__874 (
            .O(N__4201),
            .I(N__4164));
    InMux I__873 (
            .O(N__4198),
            .I(N__4164));
    InMux I__872 (
            .O(N__4197),
            .I(N__4157));
    InMux I__871 (
            .O(N__4194),
            .I(N__4157));
    InMux I__870 (
            .O(N__4191),
            .I(N__4157));
    InMux I__869 (
            .O(N__4190),
            .I(N__4146));
    InMux I__868 (
            .O(N__4189),
            .I(N__4146));
    InMux I__867 (
            .O(N__4186),
            .I(N__4146));
    InMux I__866 (
            .O(N__4183),
            .I(N__4146));
    InMux I__865 (
            .O(N__4180),
            .I(N__4146));
    InMux I__864 (
            .O(N__4177),
            .I(N__4140));
    LocalMux I__863 (
            .O(N__4164),
            .I(N__4133));
    LocalMux I__862 (
            .O(N__4157),
            .I(N__4133));
    LocalMux I__861 (
            .O(N__4146),
            .I(N__4133));
    CascadeMux I__860 (
            .O(N__4145),
            .I(N__4129));
    CascadeMux I__859 (
            .O(N__4144),
            .I(N__4125));
    CascadeMux I__858 (
            .O(N__4143),
            .I(N__4121));
    LocalMux I__857 (
            .O(N__4140),
            .I(N__4108));
    Span4Mux_v I__856 (
            .O(N__4133),
            .I(N__4105));
    InMux I__855 (
            .O(N__4132),
            .I(N__4090));
    InMux I__854 (
            .O(N__4129),
            .I(N__4090));
    InMux I__853 (
            .O(N__4128),
            .I(N__4090));
    InMux I__852 (
            .O(N__4125),
            .I(N__4090));
    InMux I__851 (
            .O(N__4124),
            .I(N__4090));
    InMux I__850 (
            .O(N__4121),
            .I(N__4090));
    InMux I__849 (
            .O(N__4120),
            .I(N__4090));
    InMux I__848 (
            .O(N__4119),
            .I(N__4087));
    CascadeMux I__847 (
            .O(N__4118),
            .I(N__4084));
    CascadeMux I__846 (
            .O(N__4117),
            .I(N__4081));
    CascadeMux I__845 (
            .O(N__4116),
            .I(N__4078));
    CascadeMux I__844 (
            .O(N__4115),
            .I(N__4075));
    CascadeMux I__843 (
            .O(N__4114),
            .I(N__4072));
    CascadeMux I__842 (
            .O(N__4113),
            .I(N__4069));
    CascadeMux I__841 (
            .O(N__4112),
            .I(N__4066));
    CascadeMux I__840 (
            .O(N__4111),
            .I(N__4063));
    Span4Mux_v I__839 (
            .O(N__4108),
            .I(N__4059));
    Span4Mux_h I__838 (
            .O(N__4105),
            .I(N__4054));
    LocalMux I__837 (
            .O(N__4090),
            .I(N__4054));
    LocalMux I__836 (
            .O(N__4087),
            .I(N__4051));
    InMux I__835 (
            .O(N__4084),
            .I(N__4042));
    InMux I__834 (
            .O(N__4081),
            .I(N__4042));
    InMux I__833 (
            .O(N__4078),
            .I(N__4042));
    InMux I__832 (
            .O(N__4075),
            .I(N__4042));
    InMux I__831 (
            .O(N__4072),
            .I(N__4033));
    InMux I__830 (
            .O(N__4069),
            .I(N__4033));
    InMux I__829 (
            .O(N__4066),
            .I(N__4033));
    InMux I__828 (
            .O(N__4063),
            .I(N__4033));
    InMux I__827 (
            .O(N__4062),
            .I(N__4030));
    Odrv4 I__826 (
            .O(N__4059),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__825 (
            .O(N__4054),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__824 (
            .O(N__4051),
            .I(CONSTANT_ONE_NET));
    LocalMux I__823 (
            .O(N__4042),
            .I(CONSTANT_ONE_NET));
    LocalMux I__822 (
            .O(N__4033),
            .I(CONSTANT_ONE_NET));
    LocalMux I__821 (
            .O(N__4030),
            .I(CONSTANT_ONE_NET));
    InMux I__820 (
            .O(N__4017),
            .I(bfn_6_9_0_));
    InMux I__819 (
            .O(N__4014),
            .I(N__4011));
    LocalMux I__818 (
            .O(N__4011),
            .I(sr_row_data_8));
    InMux I__817 (
            .O(N__4008),
            .I(N__4005));
    LocalMux I__816 (
            .O(N__4005),
            .I(N__4002));
    Odrv4 I__815 (
            .O(N__4002),
            .I(sr_row_data_6));
    InMux I__814 (
            .O(N__3999),
            .I(N__3996));
    LocalMux I__813 (
            .O(N__3996),
            .I(sr_row_data_9));
    InMux I__812 (
            .O(N__3993),
            .I(N__3990));
    LocalMux I__811 (
            .O(N__3990),
            .I(N__3987));
    Odrv4 I__810 (
            .O(N__3987),
            .I(n4));
    InMux I__809 (
            .O(N__3984),
            .I(N__3981));
    LocalMux I__808 (
            .O(N__3981),
            .I(N__3978));
    Odrv4 I__807 (
            .O(N__3978),
            .I(n5));
    InMux I__806 (
            .O(N__3975),
            .I(N__3972));
    LocalMux I__805 (
            .O(N__3972),
            .I(N__3969));
    Odrv4 I__804 (
            .O(N__3969),
            .I(n1));
    InMux I__803 (
            .O(N__3966),
            .I(N__3963));
    LocalMux I__802 (
            .O(N__3963),
            .I(n9_adj_123));
    CascadeMux I__801 (
            .O(N__3960),
            .I(n811_cascade_));
    InMux I__800 (
            .O(N__3957),
            .I(N__3954));
    LocalMux I__799 (
            .O(N__3954),
            .I(N__3951));
    Odrv4 I__798 (
            .O(N__3951),
            .I(n6));
    InMux I__797 (
            .O(N__3948),
            .I(N__3945));
    LocalMux I__796 (
            .O(N__3945),
            .I(N__3942));
    Odrv4 I__795 (
            .O(N__3942),
            .I(n12_adj_126));
    InMux I__794 (
            .O(N__3939),
            .I(N__3936));
    LocalMux I__793 (
            .O(N__3936),
            .I(n16_adj_129));
    CascadeMux I__792 (
            .O(N__3933),
            .I(n831_cascade_));
    InMux I__791 (
            .O(N__3930),
            .I(N__3927));
    LocalMux I__790 (
            .O(N__3927),
            .I(n775));
    SRMux I__789 (
            .O(N__3924),
            .I(N__3920));
    SRMux I__788 (
            .O(N__3923),
            .I(N__3916));
    LocalMux I__787 (
            .O(N__3920),
            .I(N__3910));
    SRMux I__786 (
            .O(N__3919),
            .I(N__3907));
    LocalMux I__785 (
            .O(N__3916),
            .I(N__3904));
    SRMux I__784 (
            .O(N__3915),
            .I(N__3901));
    InMux I__783 (
            .O(N__3914),
            .I(N__3898));
    InMux I__782 (
            .O(N__3913),
            .I(N__3895));
    Span4Mux_h I__781 (
            .O(N__3910),
            .I(N__3886));
    LocalMux I__780 (
            .O(N__3907),
            .I(N__3886));
    Span4Mux_h I__779 (
            .O(N__3904),
            .I(N__3881));
    LocalMux I__778 (
            .O(N__3901),
            .I(N__3881));
    LocalMux I__777 (
            .O(N__3898),
            .I(N__3872));
    LocalMux I__776 (
            .O(N__3895),
            .I(N__3872));
    InMux I__775 (
            .O(N__3894),
            .I(N__3867));
    InMux I__774 (
            .O(N__3893),
            .I(N__3867));
    InMux I__773 (
            .O(N__3892),
            .I(N__3862));
    InMux I__772 (
            .O(N__3891),
            .I(N__3862));
    Span4Mux_h I__771 (
            .O(N__3886),
            .I(N__3859));
    Span4Mux_h I__770 (
            .O(N__3881),
            .I(N__3856));
    InMux I__769 (
            .O(N__3880),
            .I(N__3851));
    InMux I__768 (
            .O(N__3879),
            .I(N__3851));
    InMux I__767 (
            .O(N__3878),
            .I(N__3846));
    InMux I__766 (
            .O(N__3877),
            .I(N__3846));
    Odrv12 I__765 (
            .O(N__3872),
            .I(reset_signal));
    LocalMux I__764 (
            .O(N__3867),
            .I(reset_signal));
    LocalMux I__763 (
            .O(N__3862),
            .I(reset_signal));
    Odrv4 I__762 (
            .O(N__3859),
            .I(reset_signal));
    Odrv4 I__761 (
            .O(N__3856),
            .I(reset_signal));
    LocalMux I__760 (
            .O(N__3851),
            .I(reset_signal));
    LocalMux I__759 (
            .O(N__3846),
            .I(reset_signal));
    CascadeMux I__758 (
            .O(N__3831),
            .I(n835_cascade_));
    InMux I__757 (
            .O(N__3828),
            .I(N__3825));
    LocalMux I__756 (
            .O(N__3825),
            .I(N__3822));
    Span4Mux_h I__755 (
            .O(N__3822),
            .I(N__3817));
    InMux I__754 (
            .O(N__3821),
            .I(N__3814));
    InMux I__753 (
            .O(N__3820),
            .I(N__3811));
    Odrv4 I__752 (
            .O(N__3817),
            .I(row_complete));
    LocalMux I__751 (
            .O(N__3814),
            .I(row_complete));
    LocalMux I__750 (
            .O(N__3811),
            .I(row_complete));
    ClkMux I__749 (
            .O(N__3804),
            .I(N__3799));
    ClkMux I__748 (
            .O(N__3803),
            .I(N__3796));
    ClkMux I__747 (
            .O(N__3802),
            .I(N__3793));
    LocalMux I__746 (
            .O(N__3799),
            .I(N__3790));
    LocalMux I__745 (
            .O(N__3796),
            .I(N__3786));
    LocalMux I__744 (
            .O(N__3793),
            .I(N__3783));
    Span4Mux_v I__743 (
            .O(N__3790),
            .I(N__3780));
    IoInMux I__742 (
            .O(N__3789),
            .I(N__3777));
    Span4Mux_h I__741 (
            .O(N__3786),
            .I(N__3774));
    Span4Mux_h I__740 (
            .O(N__3783),
            .I(N__3771));
    Span4Mux_h I__739 (
            .O(N__3780),
            .I(N__3768));
    LocalMux I__738 (
            .O(N__3777),
            .I(N__3765));
    Odrv4 I__737 (
            .O(N__3774),
            .I(divided_pulse_c));
    Odrv4 I__736 (
            .O(N__3771),
            .I(divided_pulse_c));
    Odrv4 I__735 (
            .O(N__3768),
            .I(divided_pulse_c));
    Odrv12 I__734 (
            .O(N__3765),
            .I(divided_pulse_c));
    InMux I__733 (
            .O(N__3756),
            .I(N__3752));
    InMux I__732 (
            .O(N__3755),
            .I(N__3749));
    LocalMux I__731 (
            .O(N__3752),
            .I(\row_counter.internal_count_8 ));
    LocalMux I__730 (
            .O(N__3749),
            .I(\row_counter.internal_count_8 ));
    InMux I__729 (
            .O(N__3744),
            .I(bfn_6_8_0_));
    InMux I__728 (
            .O(N__3741),
            .I(N__3737));
    InMux I__727 (
            .O(N__3740),
            .I(N__3734));
    LocalMux I__726 (
            .O(N__3737),
            .I(N__3731));
    LocalMux I__725 (
            .O(N__3734),
            .I(\row_counter.internal_count_9 ));
    Odrv4 I__724 (
            .O(N__3731),
            .I(\row_counter.internal_count_9 ));
    InMux I__723 (
            .O(N__3726),
            .I(\row_counter.n704 ));
    InMux I__722 (
            .O(N__3723),
            .I(N__3719));
    InMux I__721 (
            .O(N__3722),
            .I(N__3716));
    LocalMux I__720 (
            .O(N__3719),
            .I(\row_counter.internal_count_10 ));
    LocalMux I__719 (
            .O(N__3716),
            .I(\row_counter.internal_count_10 ));
    InMux I__718 (
            .O(N__3711),
            .I(\row_counter.n705 ));
    InMux I__717 (
            .O(N__3708),
            .I(N__3704));
    InMux I__716 (
            .O(N__3707),
            .I(N__3701));
    LocalMux I__715 (
            .O(N__3704),
            .I(\row_counter.internal_count_11 ));
    LocalMux I__714 (
            .O(N__3701),
            .I(\row_counter.internal_count_11 ));
    InMux I__713 (
            .O(N__3696),
            .I(\row_counter.n706 ));
    InMux I__712 (
            .O(N__3693),
            .I(N__3689));
    InMux I__711 (
            .O(N__3692),
            .I(N__3686));
    LocalMux I__710 (
            .O(N__3689),
            .I(\row_counter.internal_count_12 ));
    LocalMux I__709 (
            .O(N__3686),
            .I(\row_counter.internal_count_12 ));
    InMux I__708 (
            .O(N__3681),
            .I(\row_counter.n707 ));
    InMux I__707 (
            .O(N__3678),
            .I(N__3674));
    InMux I__706 (
            .O(N__3677),
            .I(N__3671));
    LocalMux I__705 (
            .O(N__3674),
            .I(\row_counter.internal_count_13 ));
    LocalMux I__704 (
            .O(N__3671),
            .I(\row_counter.internal_count_13 ));
    InMux I__703 (
            .O(N__3666),
            .I(\row_counter.n708 ));
    InMux I__702 (
            .O(N__3663),
            .I(N__3659));
    InMux I__701 (
            .O(N__3662),
            .I(N__3656));
    LocalMux I__700 (
            .O(N__3659),
            .I(\row_counter.internal_count_14 ));
    LocalMux I__699 (
            .O(N__3656),
            .I(\row_counter.internal_count_14 ));
    InMux I__698 (
            .O(N__3651),
            .I(\row_counter.n709 ));
    InMux I__697 (
            .O(N__3648),
            .I(N__3644));
    InMux I__696 (
            .O(N__3647),
            .I(N__3641));
    LocalMux I__695 (
            .O(N__3644),
            .I(\row_counter.internal_count_15 ));
    LocalMux I__694 (
            .O(N__3641),
            .I(\row_counter.internal_count_15 ));
    InMux I__693 (
            .O(N__3636),
            .I(\row_counter.n710 ));
    InMux I__692 (
            .O(N__3633),
            .I(N__3624));
    InMux I__691 (
            .O(N__3632),
            .I(N__3624));
    InMux I__690 (
            .O(N__3631),
            .I(N__3624));
    LocalMux I__689 (
            .O(N__3624),
            .I(shifted_data_1_adj_114));
    InMux I__688 (
            .O(N__3621),
            .I(N__3617));
    InMux I__687 (
            .O(N__3620),
            .I(N__3614));
    LocalMux I__686 (
            .O(N__3617),
            .I(\row_counter.internal_count_0 ));
    LocalMux I__685 (
            .O(N__3614),
            .I(\row_counter.internal_count_0 ));
    InMux I__684 (
            .O(N__3609),
            .I(N__3606));
    LocalMux I__683 (
            .O(N__3606),
            .I(N__3603));
    Odrv4 I__682 (
            .O(N__3603),
            .I(sr_row_data_0));
    InMux I__681 (
            .O(N__3600),
            .I(bfn_6_7_0_));
    InMux I__680 (
            .O(N__3597),
            .I(N__3593));
    InMux I__679 (
            .O(N__3596),
            .I(N__3590));
    LocalMux I__678 (
            .O(N__3593),
            .I(\row_counter.internal_count_1 ));
    LocalMux I__677 (
            .O(N__3590),
            .I(\row_counter.internal_count_1 ));
    CascadeMux I__676 (
            .O(N__3585),
            .I(N__3582));
    InMux I__675 (
            .O(N__3582),
            .I(N__3579));
    LocalMux I__674 (
            .O(N__3579),
            .I(sr_row_data_1));
    InMux I__673 (
            .O(N__3576),
            .I(\row_counter.n696 ));
    InMux I__672 (
            .O(N__3573),
            .I(N__3569));
    InMux I__671 (
            .O(N__3572),
            .I(N__3566));
    LocalMux I__670 (
            .O(N__3569),
            .I(N__3561));
    LocalMux I__669 (
            .O(N__3566),
            .I(N__3561));
    Odrv4 I__668 (
            .O(N__3561),
            .I(\row_counter.internal_count_2 ));
    InMux I__667 (
            .O(N__3558),
            .I(\row_counter.n697 ));
    InMux I__666 (
            .O(N__3555),
            .I(N__3552));
    LocalMux I__665 (
            .O(N__3552),
            .I(N__3548));
    InMux I__664 (
            .O(N__3551),
            .I(N__3545));
    Odrv4 I__663 (
            .O(N__3548),
            .I(\row_counter.internal_count_3 ));
    LocalMux I__662 (
            .O(N__3545),
            .I(\row_counter.internal_count_3 ));
    InMux I__661 (
            .O(N__3540),
            .I(\row_counter.n698 ));
    InMux I__660 (
            .O(N__3537),
            .I(N__3533));
    InMux I__659 (
            .O(N__3536),
            .I(N__3530));
    LocalMux I__658 (
            .O(N__3533),
            .I(\row_counter.internal_count_4 ));
    LocalMux I__657 (
            .O(N__3530),
            .I(\row_counter.internal_count_4 ));
    InMux I__656 (
            .O(N__3525),
            .I(N__3522));
    LocalMux I__655 (
            .O(N__3522),
            .I(N__3519));
    Odrv4 I__654 (
            .O(N__3519),
            .I(sr_row_data_4));
    InMux I__653 (
            .O(N__3516),
            .I(\row_counter.n699 ));
    InMux I__652 (
            .O(N__3513),
            .I(N__3509));
    InMux I__651 (
            .O(N__3512),
            .I(N__3506));
    LocalMux I__650 (
            .O(N__3509),
            .I(\row_counter.internal_count_5 ));
    LocalMux I__649 (
            .O(N__3506),
            .I(\row_counter.internal_count_5 ));
    InMux I__648 (
            .O(N__3501),
            .I(\row_counter.n700 ));
    InMux I__647 (
            .O(N__3498),
            .I(N__3494));
    InMux I__646 (
            .O(N__3497),
            .I(N__3491));
    LocalMux I__645 (
            .O(N__3494),
            .I(\row_counter.internal_count_6 ));
    LocalMux I__644 (
            .O(N__3491),
            .I(\row_counter.internal_count_6 ));
    InMux I__643 (
            .O(N__3486),
            .I(\row_counter.n701 ));
    InMux I__642 (
            .O(N__3483),
            .I(N__3479));
    InMux I__641 (
            .O(N__3482),
            .I(N__3476));
    LocalMux I__640 (
            .O(N__3479),
            .I(\row_counter.internal_count_7 ));
    LocalMux I__639 (
            .O(N__3476),
            .I(\row_counter.internal_count_7 ));
    CascadeMux I__638 (
            .O(N__3471),
            .I(N__3468));
    InMux I__637 (
            .O(N__3468),
            .I(N__3465));
    LocalMux I__636 (
            .O(N__3465),
            .I(N__3462));
    Odrv4 I__635 (
            .O(N__3462),
            .I(sr_row_data_7));
    InMux I__634 (
            .O(N__3459),
            .I(\row_counter.n702 ));
    InMux I__633 (
            .O(N__3456),
            .I(N__3453));
    LocalMux I__632 (
            .O(N__3453),
            .I(N__3450));
    Span4Mux_h I__631 (
            .O(N__3450),
            .I(N__3447));
    Sp12to4 I__630 (
            .O(N__3447),
            .I(N__3444));
    Span12Mux_v I__629 (
            .O(N__3444),
            .I(N__3441));
    Odrv12 I__628 (
            .O(N__3441),
            .I(en_rowpack_c));
    CEMux I__627 (
            .O(N__3438),
            .I(N__3434));
    CEMux I__626 (
            .O(N__3437),
            .I(N__3431));
    LocalMux I__625 (
            .O(N__3434),
            .I(N__3428));
    LocalMux I__624 (
            .O(N__3431),
            .I(N__3425));
    Odrv12 I__623 (
            .O(N__3428),
            .I(n189));
    Odrv4 I__622 (
            .O(N__3425),
            .I(n189));
    InMux I__621 (
            .O(N__3420),
            .I(N__3417));
    LocalMux I__620 (
            .O(N__3417),
            .I(N__3413));
    InMux I__619 (
            .O(N__3416),
            .I(N__3410));
    Span4Mux_v I__618 (
            .O(N__3413),
            .I(N__3405));
    LocalMux I__617 (
            .O(N__3410),
            .I(N__3405));
    Span4Mux_v I__616 (
            .O(N__3405),
            .I(N__3402));
    Span4Mux_v I__615 (
            .O(N__3402),
            .I(N__3399));
    Sp12to4 I__614 (
            .O(N__3399),
            .I(N__3396));
    Odrv12 I__613 (
            .O(N__3396),
            .I(sr_data_c));
    InMux I__612 (
            .O(N__3393),
            .I(N__3390));
    LocalMux I__611 (
            .O(N__3390),
            .I(N__3385));
    InMux I__610 (
            .O(N__3389),
            .I(N__3380));
    InMux I__609 (
            .O(N__3388),
            .I(N__3380));
    Odrv4 I__608 (
            .O(N__3385),
            .I(shifted_data_0));
    LocalMux I__607 (
            .O(N__3380),
            .I(shifted_data_0));
    InMux I__606 (
            .O(N__3375),
            .I(N__3371));
    CascadeMux I__605 (
            .O(N__3374),
            .I(N__3368));
    LocalMux I__604 (
            .O(N__3371),
            .I(N__3364));
    InMux I__603 (
            .O(N__3368),
            .I(N__3361));
    InMux I__602 (
            .O(N__3367),
            .I(N__3358));
    Odrv4 I__601 (
            .O(N__3364),
            .I(shifted_data_1));
    LocalMux I__600 (
            .O(N__3361),
            .I(shifted_data_1));
    LocalMux I__599 (
            .O(N__3358),
            .I(shifted_data_1));
    CascadeMux I__598 (
            .O(N__3351),
            .I(N__3347));
    InMux I__597 (
            .O(N__3350),
            .I(N__3344));
    InMux I__596 (
            .O(N__3347),
            .I(N__3340));
    LocalMux I__595 (
            .O(N__3344),
            .I(N__3337));
    InMux I__594 (
            .O(N__3343),
            .I(N__3334));
    LocalMux I__593 (
            .O(N__3340),
            .I(N__3331));
    Odrv12 I__592 (
            .O(N__3337),
            .I(shifted_data_2));
    LocalMux I__591 (
            .O(N__3334),
            .I(shifted_data_2));
    Odrv4 I__590 (
            .O(N__3331),
            .I(shifted_data_2));
    InMux I__589 (
            .O(N__3324),
            .I(N__3321));
    LocalMux I__588 (
            .O(N__3321),
            .I(N__3312));
    InMux I__587 (
            .O(N__3320),
            .I(N__3303));
    InMux I__586 (
            .O(N__3319),
            .I(N__3303));
    InMux I__585 (
            .O(N__3318),
            .I(N__3303));
    InMux I__584 (
            .O(N__3317),
            .I(N__3303));
    CascadeMux I__583 (
            .O(N__3316),
            .I(N__3299));
    CascadeMux I__582 (
            .O(N__3315),
            .I(N__3291));
    Span4Mux_v I__581 (
            .O(N__3312),
            .I(N__3286));
    LocalMux I__580 (
            .O(N__3303),
            .I(N__3283));
    InMux I__579 (
            .O(N__3302),
            .I(N__3270));
    InMux I__578 (
            .O(N__3299),
            .I(N__3270));
    InMux I__577 (
            .O(N__3298),
            .I(N__3270));
    InMux I__576 (
            .O(N__3297),
            .I(N__3270));
    InMux I__575 (
            .O(N__3296),
            .I(N__3270));
    InMux I__574 (
            .O(N__3295),
            .I(N__3270));
    InMux I__573 (
            .O(N__3294),
            .I(N__3261));
    InMux I__572 (
            .O(N__3291),
            .I(N__3261));
    InMux I__571 (
            .O(N__3290),
            .I(N__3261));
    InMux I__570 (
            .O(N__3289),
            .I(N__3261));
    Odrv4 I__569 (
            .O(N__3286),
            .I(n330));
    Odrv12 I__568 (
            .O(N__3283),
            .I(n330));
    LocalMux I__567 (
            .O(N__3270),
            .I(n330));
    LocalMux I__566 (
            .O(N__3261),
            .I(n330));
    CascadeMux I__565 (
            .O(N__3252),
            .I(N__3249));
    InMux I__564 (
            .O(N__3249),
            .I(N__3245));
    CascadeMux I__563 (
            .O(N__3248),
            .I(N__3239));
    LocalMux I__562 (
            .O(N__3245),
            .I(N__3233));
    InMux I__561 (
            .O(N__3244),
            .I(N__3228));
    InMux I__560 (
            .O(N__3243),
            .I(N__3228));
    InMux I__559 (
            .O(N__3242),
            .I(N__3223));
    InMux I__558 (
            .O(N__3239),
            .I(N__3223));
    CascadeMux I__557 (
            .O(N__3238),
            .I(N__3217));
    CascadeMux I__556 (
            .O(N__3237),
            .I(N__3213));
    CascadeMux I__555 (
            .O(N__3236),
            .I(N__3207));
    Span4Mux_v I__554 (
            .O(N__3233),
            .I(N__3204));
    LocalMux I__553 (
            .O(N__3228),
            .I(N__3199));
    LocalMux I__552 (
            .O(N__3223),
            .I(N__3199));
    InMux I__551 (
            .O(N__3222),
            .I(N__3186));
    InMux I__550 (
            .O(N__3221),
            .I(N__3186));
    InMux I__549 (
            .O(N__3220),
            .I(N__3186));
    InMux I__548 (
            .O(N__3217),
            .I(N__3186));
    InMux I__547 (
            .O(N__3216),
            .I(N__3186));
    InMux I__546 (
            .O(N__3213),
            .I(N__3186));
    InMux I__545 (
            .O(N__3212),
            .I(N__3183));
    InMux I__544 (
            .O(N__3211),
            .I(N__3176));
    InMux I__543 (
            .O(N__3210),
            .I(N__3176));
    InMux I__542 (
            .O(N__3207),
            .I(N__3176));
    Odrv4 I__541 (
            .O(N__3204),
            .I(n169));
    Odrv12 I__540 (
            .O(N__3199),
            .I(n169));
    LocalMux I__539 (
            .O(N__3186),
            .I(n169));
    LocalMux I__538 (
            .O(N__3183),
            .I(n169));
    LocalMux I__537 (
            .O(N__3176),
            .I(n169));
    InMux I__536 (
            .O(N__3165),
            .I(N__3161));
    CascadeMux I__535 (
            .O(N__3164),
            .I(N__3157));
    LocalMux I__534 (
            .O(N__3161),
            .I(N__3154));
    InMux I__533 (
            .O(N__3160),
            .I(N__3151));
    InMux I__532 (
            .O(N__3157),
            .I(N__3148));
    Odrv4 I__531 (
            .O(N__3154),
            .I(shifted_data_3));
    LocalMux I__530 (
            .O(N__3151),
            .I(shifted_data_3));
    LocalMux I__529 (
            .O(N__3148),
            .I(shifted_data_3));
    CascadeMux I__528 (
            .O(N__3141),
            .I(N__3137));
    InMux I__527 (
            .O(N__3140),
            .I(N__3134));
    InMux I__526 (
            .O(N__3137),
            .I(N__3130));
    LocalMux I__525 (
            .O(N__3134),
            .I(N__3127));
    InMux I__524 (
            .O(N__3133),
            .I(N__3124));
    LocalMux I__523 (
            .O(N__3130),
            .I(N__3121));
    Odrv12 I__522 (
            .O(N__3127),
            .I(shifted_data_4));
    LocalMux I__521 (
            .O(N__3124),
            .I(shifted_data_4));
    Odrv4 I__520 (
            .O(N__3121),
            .I(shifted_data_4));
    InMux I__519 (
            .O(N__3114),
            .I(N__3111));
    LocalMux I__518 (
            .O(N__3111),
            .I(N__3106));
    InMux I__517 (
            .O(N__3110),
            .I(N__3103));
    InMux I__516 (
            .O(N__3109),
            .I(N__3100));
    Odrv4 I__515 (
            .O(N__3106),
            .I(shifted_data_0_adj_115));
    LocalMux I__514 (
            .O(N__3103),
            .I(shifted_data_0_adj_115));
    LocalMux I__513 (
            .O(N__3100),
            .I(shifted_data_0_adj_115));
    InMux I__512 (
            .O(N__3093),
            .I(\row_counter.n752 ));
    InMux I__511 (
            .O(N__3090),
            .I(\row_counter.n753 ));
    InMux I__510 (
            .O(N__3087),
            .I(\row_counter.n754 ));
    InMux I__509 (
            .O(N__3084),
            .I(\row_counter.n755 ));
    InMux I__508 (
            .O(N__3081),
            .I(\row_counter.n756 ));
    InMux I__507 (
            .O(N__3078),
            .I(\row_counter.n757 ));
    InMux I__506 (
            .O(N__3075),
            .I(\row_counter.n743 ));
    InMux I__505 (
            .O(N__3072),
            .I(\row_counter.n744 ));
    InMux I__504 (
            .O(N__3069),
            .I(\row_counter.n745 ));
    InMux I__503 (
            .O(N__3066),
            .I(\row_counter.n746 ));
    InMux I__502 (
            .O(N__3063),
            .I(\row_counter.n747 ));
    InMux I__501 (
            .O(N__3060),
            .I(\row_counter.n748 ));
    InMux I__500 (
            .O(N__3057),
            .I(\row_counter.n749 ));
    InMux I__499 (
            .O(N__3054),
            .I(bfn_5_8_0_));
    InMux I__498 (
            .O(N__3051),
            .I(\row_counter.n751 ));
    CascadeMux I__497 (
            .O(N__3048),
            .I(N__3044));
    InMux I__496 (
            .O(N__3047),
            .I(N__3040));
    InMux I__495 (
            .O(N__3044),
            .I(N__3037));
    InMux I__494 (
            .O(N__3043),
            .I(N__3034));
    LocalMux I__493 (
            .O(N__3040),
            .I(shifted_data_12));
    LocalMux I__492 (
            .O(N__3037),
            .I(shifted_data_12));
    LocalMux I__491 (
            .O(N__3034),
            .I(shifted_data_12));
    InMux I__490 (
            .O(N__3027),
            .I(N__3022));
    InMux I__489 (
            .O(N__3026),
            .I(N__3017));
    InMux I__488 (
            .O(N__3025),
            .I(N__3017));
    LocalMux I__487 (
            .O(N__3022),
            .I(shifted_data_13));
    LocalMux I__486 (
            .O(N__3017),
            .I(shifted_data_13));
    InMux I__485 (
            .O(N__3012),
            .I(N__3007));
    InMux I__484 (
            .O(N__3011),
            .I(N__3002));
    InMux I__483 (
            .O(N__3010),
            .I(N__3002));
    LocalMux I__482 (
            .O(N__3007),
            .I(shifted_data_8));
    LocalMux I__481 (
            .O(N__3002),
            .I(shifted_data_8));
    CascadeMux I__480 (
            .O(N__2997),
            .I(N__2993));
    InMux I__479 (
            .O(N__2996),
            .I(N__2989));
    InMux I__478 (
            .O(N__2993),
            .I(N__2986));
    InMux I__477 (
            .O(N__2992),
            .I(N__2983));
    LocalMux I__476 (
            .O(N__2989),
            .I(shifted_data_9));
    LocalMux I__475 (
            .O(N__2986),
            .I(shifted_data_9));
    LocalMux I__474 (
            .O(N__2983),
            .I(shifted_data_9));
    InMux I__473 (
            .O(N__2976),
            .I(N__2971));
    InMux I__472 (
            .O(N__2975),
            .I(N__2968));
    InMux I__471 (
            .O(N__2974),
            .I(N__2965));
    LocalMux I__470 (
            .O(N__2971),
            .I(shifted_data_10));
    LocalMux I__469 (
            .O(N__2968),
            .I(shifted_data_10));
    LocalMux I__468 (
            .O(N__2965),
            .I(shifted_data_10));
    InMux I__467 (
            .O(N__2958),
            .I(N__2953));
    InMux I__466 (
            .O(N__2957),
            .I(N__2948));
    InMux I__465 (
            .O(N__2956),
            .I(N__2948));
    LocalMux I__464 (
            .O(N__2953),
            .I(shifted_data_5));
    LocalMux I__463 (
            .O(N__2948),
            .I(shifted_data_5));
    InMux I__462 (
            .O(N__2943),
            .I(N__2938));
    InMux I__461 (
            .O(N__2942),
            .I(N__2933));
    InMux I__460 (
            .O(N__2941),
            .I(N__2933));
    LocalMux I__459 (
            .O(N__2938),
            .I(shifted_data_6));
    LocalMux I__458 (
            .O(N__2933),
            .I(shifted_data_6));
    CascadeMux I__457 (
            .O(N__2928),
            .I(N__2924));
    InMux I__456 (
            .O(N__2927),
            .I(N__2920));
    InMux I__455 (
            .O(N__2924),
            .I(N__2917));
    InMux I__454 (
            .O(N__2923),
            .I(N__2914));
    LocalMux I__453 (
            .O(N__2920),
            .I(shifted_data_7));
    LocalMux I__452 (
            .O(N__2917),
            .I(shifted_data_7));
    LocalMux I__451 (
            .O(N__2914),
            .I(shifted_data_7));
    InMux I__450 (
            .O(N__2907),
            .I(bfn_5_7_0_));
    InMux I__449 (
            .O(N__2904),
            .I(N__2901));
    LocalMux I__448 (
            .O(N__2901),
            .I(n2_adj_99));
    InMux I__447 (
            .O(N__2898),
            .I(N__2895));
    LocalMux I__446 (
            .O(N__2895),
            .I(n11));
    CascadeMux I__445 (
            .O(N__2892),
            .I(n823_cascade_));
    InMux I__444 (
            .O(N__2889),
            .I(N__2886));
    LocalMux I__443 (
            .O(N__2886),
            .I(n781));
    InMux I__442 (
            .O(N__2883),
            .I(N__2880));
    LocalMux I__441 (
            .O(N__2880),
            .I(n827));
    InMux I__440 (
            .O(N__2877),
            .I(N__2871));
    InMux I__439 (
            .O(N__2876),
            .I(N__2871));
    LocalMux I__438 (
            .O(N__2871),
            .I(N__2868));
    Span4Mux_v I__437 (
            .O(N__2868),
            .I(N__2865));
    Sp12to4 I__436 (
            .O(N__2865),
            .I(N__2862));
    Odrv12 I__435 (
            .O(N__2862),
            .I(sr_sel_row_c));
    CascadeMux I__434 (
            .O(N__2859),
            .I(n169_cascade_));
    InMux I__433 (
            .O(N__2856),
            .I(N__2850));
    InMux I__432 (
            .O(N__2855),
            .I(N__2850));
    LocalMux I__431 (
            .O(N__2850),
            .I(N__2847));
    Span12Mux_h I__430 (
            .O(N__2847),
            .I(N__2844));
    Span12Mux_v I__429 (
            .O(N__2844),
            .I(N__2841));
    Odrv12 I__428 (
            .O(N__2841),
            .I(sr_sel_div_c));
    InMux I__427 (
            .O(N__2838),
            .I(N__2830));
    InMux I__426 (
            .O(N__2837),
            .I(N__2830));
    InMux I__425 (
            .O(N__2836),
            .I(N__2825));
    InMux I__424 (
            .O(N__2835),
            .I(N__2825));
    LocalMux I__423 (
            .O(N__2830),
            .I(N__2820));
    LocalMux I__422 (
            .O(N__2825),
            .I(N__2820));
    Span4Mux_v I__421 (
            .O(N__2820),
            .I(N__2817));
    Sp12to4 I__420 (
            .O(N__2817),
            .I(N__2814));
    Odrv12 I__419 (
            .O(N__2814),
            .I(sr_reset_c));
    CascadeMux I__418 (
            .O(N__2811),
            .I(n330_cascade_));
    InMux I__417 (
            .O(N__2808),
            .I(N__2803));
    InMux I__416 (
            .O(N__2807),
            .I(N__2798));
    InMux I__415 (
            .O(N__2806),
            .I(N__2798));
    LocalMux I__414 (
            .O(N__2803),
            .I(shifted_data_14));
    LocalMux I__413 (
            .O(N__2798),
            .I(shifted_data_14));
    InMux I__412 (
            .O(N__2793),
            .I(N__2789));
    InMux I__411 (
            .O(N__2792),
            .I(N__2786));
    LocalMux I__410 (
            .O(N__2789),
            .I(shifted_data_15));
    LocalMux I__409 (
            .O(N__2786),
            .I(shifted_data_15));
    InMux I__408 (
            .O(N__2781),
            .I(N__2776));
    InMux I__407 (
            .O(N__2780),
            .I(N__2771));
    InMux I__406 (
            .O(N__2779),
            .I(N__2771));
    LocalMux I__405 (
            .O(N__2776),
            .I(shifted_data_11));
    LocalMux I__404 (
            .O(N__2771),
            .I(shifted_data_11));
    InMux I__403 (
            .O(N__2766),
            .I(N__2763));
    LocalMux I__402 (
            .O(N__2763),
            .I(N__2760));
    Odrv4 I__401 (
            .O(N__2760),
            .I(sr_divider_data_10));
    InMux I__400 (
            .O(N__2757),
            .I(N__2754));
    LocalMux I__399 (
            .O(N__2754),
            .I(N__2751));
    Odrv12 I__398 (
            .O(N__2751),
            .I(sr_divider_data_6));
    InMux I__397 (
            .O(N__2748),
            .I(N__2745));
    LocalMux I__396 (
            .O(N__2745),
            .I(N__2742));
    Odrv4 I__395 (
            .O(N__2742),
            .I(sr_divider_data_9));
    CascadeMux I__394 (
            .O(N__2739),
            .I(N__2736));
    InMux I__393 (
            .O(N__2736),
            .I(N__2733));
    LocalMux I__392 (
            .O(N__2733),
            .I(N__2730));
    Odrv12 I__391 (
            .O(N__2730),
            .I(sr_divider_data_4));
    InMux I__390 (
            .O(N__2727),
            .I(N__2724));
    LocalMux I__389 (
            .O(N__2724),
            .I(N__2721));
    Odrv12 I__388 (
            .O(N__2721),
            .I(sr_divider_data_5));
    InMux I__387 (
            .O(N__2718),
            .I(N__2715));
    LocalMux I__386 (
            .O(N__2715),
            .I(N__2712));
    Span4Mux_v I__385 (
            .O(N__2712),
            .I(N__2709));
    Odrv4 I__384 (
            .O(N__2709),
            .I(sr_divider_data_8));
    InMux I__383 (
            .O(N__2706),
            .I(N__2703));
    LocalMux I__382 (
            .O(N__2703),
            .I(N__2700));
    Odrv12 I__381 (
            .O(N__2700),
            .I(sr_divider_data_7));
    InMux I__380 (
            .O(N__2697),
            .I(N__2694));
    LocalMux I__379 (
            .O(N__2694),
            .I(n8));
    InMux I__378 (
            .O(N__2691),
            .I(N__2688));
    LocalMux I__377 (
            .O(N__2688),
            .I(n3_adj_118));
    InMux I__376 (
            .O(N__2685),
            .I(N__2682));
    LocalMux I__375 (
            .O(N__2682),
            .I(n15));
    InMux I__374 (
            .O(N__2679),
            .I(N__2676));
    LocalMux I__373 (
            .O(N__2676),
            .I(n7));
    CascadeMux I__372 (
            .O(N__2673),
            .I(N__2670));
    InMux I__371 (
            .O(N__2670),
            .I(N__2667));
    LocalMux I__370 (
            .O(N__2667),
            .I(n10));
    InMux I__369 (
            .O(N__2664),
            .I(N__2661));
    LocalMux I__368 (
            .O(N__2661),
            .I(n14));
    CascadeMux I__367 (
            .O(N__2658),
            .I(N__2655));
    InMux I__366 (
            .O(N__2655),
            .I(N__2652));
    LocalMux I__365 (
            .O(N__2652),
            .I(sr_divider_data_13));
    InMux I__364 (
            .O(N__2649),
            .I(N__2641));
    InMux I__363 (
            .O(N__2648),
            .I(N__2641));
    InMux I__362 (
            .O(N__2647),
            .I(N__2636));
    InMux I__361 (
            .O(N__2646),
            .I(N__2636));
    LocalMux I__360 (
            .O(N__2641),
            .I(count_done));
    LocalMux I__359 (
            .O(N__2636),
            .I(count_done));
    ClkMux I__358 (
            .O(N__2631),
            .I(N__2619));
    ClkMux I__357 (
            .O(N__2630),
            .I(N__2619));
    ClkMux I__356 (
            .O(N__2629),
            .I(N__2619));
    ClkMux I__355 (
            .O(N__2628),
            .I(N__2619));
    GlobalMux I__354 (
            .O(N__2619),
            .I(N__2616));
    gio2CtrlBuf I__353 (
            .O(N__2616),
            .I(laser_pulse_c));
    CascadeMux I__352 (
            .O(N__2613),
            .I(N__2610));
    InMux I__351 (
            .O(N__2610),
            .I(N__2607));
    LocalMux I__350 (
            .O(N__2607),
            .I(N__2604));
    Odrv12 I__349 (
            .O(N__2604),
            .I(sr_divider_data_2));
    CascadeMux I__348 (
            .O(N__2601),
            .I(N__2598));
    InMux I__347 (
            .O(N__2598),
            .I(N__2595));
    LocalMux I__346 (
            .O(N__2595),
            .I(N__2592));
    Odrv12 I__345 (
            .O(N__2592),
            .I(sr_divider_data_14));
    CascadeMux I__344 (
            .O(N__2589),
            .I(N__2586));
    InMux I__343 (
            .O(N__2586),
            .I(N__2583));
    LocalMux I__342 (
            .O(N__2583),
            .I(N__2580));
    Odrv4 I__341 (
            .O(N__2580),
            .I(sr_divider_data_15));
    InMux I__340 (
            .O(N__2577),
            .I(N__2574));
    LocalMux I__339 (
            .O(N__2574),
            .I(N__2571));
    Odrv4 I__338 (
            .O(N__2571),
            .I(sr_divider_data_0));
    InMux I__337 (
            .O(N__2568),
            .I(N__2565));
    LocalMux I__336 (
            .O(N__2565),
            .I(N__2562));
    Odrv4 I__335 (
            .O(N__2562),
            .I(sr_divider_data_3));
    InMux I__334 (
            .O(N__2559),
            .I(N__2556));
    LocalMux I__333 (
            .O(N__2556),
            .I(N__2553));
    Odrv4 I__332 (
            .O(N__2553),
            .I(sr_divider_data_12));
    InMux I__331 (
            .O(N__2550),
            .I(N__2547));
    LocalMux I__330 (
            .O(N__2547),
            .I(N__2544));
    Odrv12 I__329 (
            .O(N__2544),
            .I(sr_divider_data_1));
    InMux I__328 (
            .O(N__2541),
            .I(N__2537));
    InMux I__327 (
            .O(N__2540),
            .I(N__2534));
    LocalMux I__326 (
            .O(N__2537),
            .I(N__2531));
    LocalMux I__325 (
            .O(N__2534),
            .I(\pulse_counter.internal_count_14 ));
    Odrv4 I__324 (
            .O(N__2531),
            .I(\pulse_counter.internal_count_14 ));
    InMux I__323 (
            .O(N__2526),
            .I(\pulse_counter.n725 ));
    InMux I__322 (
            .O(N__2523),
            .I(N__2519));
    InMux I__321 (
            .O(N__2522),
            .I(N__2516));
    LocalMux I__320 (
            .O(N__2519),
            .I(N__2513));
    LocalMux I__319 (
            .O(N__2516),
            .I(\pulse_counter.internal_count_15 ));
    Odrv4 I__318 (
            .O(N__2513),
            .I(\pulse_counter.internal_count_15 ));
    InMux I__317 (
            .O(N__2508),
            .I(\pulse_counter.n726 ));
    InMux I__316 (
            .O(N__2505),
            .I(N__2502));
    LocalMux I__315 (
            .O(N__2502),
            .I(\pulse_counter.n13 ));
    InMux I__314 (
            .O(N__2499),
            .I(bfn_2_9_0_));
    InMux I__313 (
            .O(N__2496),
            .I(N__2493));
    LocalMux I__312 (
            .O(N__2493),
            .I(N__2490));
    Odrv4 I__311 (
            .O(N__2490),
            .I(n4_adj_116));
    InMux I__310 (
            .O(N__2487),
            .I(N__2484));
    LocalMux I__309 (
            .O(N__2484),
            .I(N__2481));
    Odrv4 I__308 (
            .O(N__2481),
            .I(n5_adj_120));
    InMux I__307 (
            .O(N__2478),
            .I(N__2475));
    LocalMux I__306 (
            .O(N__2475),
            .I(N__2472));
    Odrv4 I__305 (
            .O(N__2472),
            .I(n1_adj_117));
    InMux I__304 (
            .O(N__2469),
            .I(N__2466));
    LocalMux I__303 (
            .O(N__2466),
            .I(n9));
    CascadeMux I__302 (
            .O(N__2463),
            .I(n795_cascade_));
    InMux I__301 (
            .O(N__2460),
            .I(N__2457));
    LocalMux I__300 (
            .O(N__2457),
            .I(N__2454));
    Odrv4 I__299 (
            .O(N__2454),
            .I(n6_adj_119));
    InMux I__298 (
            .O(N__2451),
            .I(N__2448));
    LocalMux I__297 (
            .O(N__2448),
            .I(n12));
    InMux I__296 (
            .O(N__2445),
            .I(N__2442));
    LocalMux I__295 (
            .O(N__2442),
            .I(n16));
    CascadeMux I__294 (
            .O(N__2439),
            .I(n817_cascade_));
    InMux I__293 (
            .O(N__2436),
            .I(N__2433));
    LocalMux I__292 (
            .O(N__2433),
            .I(n787));
    CascadeMux I__291 (
            .O(N__2430),
            .I(n825_cascade_));
    InMux I__290 (
            .O(N__2427),
            .I(N__2424));
    LocalMux I__289 (
            .O(N__2424),
            .I(sr_divider_data_11));
    InMux I__288 (
            .O(N__2421),
            .I(N__2417));
    InMux I__287 (
            .O(N__2420),
            .I(N__2414));
    LocalMux I__286 (
            .O(N__2417),
            .I(\pulse_counter.internal_count_5 ));
    LocalMux I__285 (
            .O(N__2414),
            .I(\pulse_counter.internal_count_5 ));
    InMux I__284 (
            .O(N__2409),
            .I(\pulse_counter.n716 ));
    InMux I__283 (
            .O(N__2406),
            .I(N__2402));
    InMux I__282 (
            .O(N__2405),
            .I(N__2399));
    LocalMux I__281 (
            .O(N__2402),
            .I(\pulse_counter.internal_count_6 ));
    LocalMux I__280 (
            .O(N__2399),
            .I(\pulse_counter.internal_count_6 ));
    InMux I__279 (
            .O(N__2394),
            .I(\pulse_counter.n717 ));
    InMux I__278 (
            .O(N__2391),
            .I(N__2387));
    InMux I__277 (
            .O(N__2390),
            .I(N__2384));
    LocalMux I__276 (
            .O(N__2387),
            .I(\pulse_counter.internal_count_7 ));
    LocalMux I__275 (
            .O(N__2384),
            .I(\pulse_counter.internal_count_7 ));
    InMux I__274 (
            .O(N__2379),
            .I(\pulse_counter.n718 ));
    InMux I__273 (
            .O(N__2376),
            .I(N__2372));
    InMux I__272 (
            .O(N__2375),
            .I(N__2369));
    LocalMux I__271 (
            .O(N__2372),
            .I(\pulse_counter.internal_count_8 ));
    LocalMux I__270 (
            .O(N__2369),
            .I(\pulse_counter.internal_count_8 ));
    InMux I__269 (
            .O(N__2364),
            .I(bfn_2_8_0_));
    InMux I__268 (
            .O(N__2361),
            .I(N__2357));
    InMux I__267 (
            .O(N__2360),
            .I(N__2354));
    LocalMux I__266 (
            .O(N__2357),
            .I(\pulse_counter.internal_count_9 ));
    LocalMux I__265 (
            .O(N__2354),
            .I(\pulse_counter.internal_count_9 ));
    InMux I__264 (
            .O(N__2349),
            .I(\pulse_counter.n720 ));
    InMux I__263 (
            .O(N__2346),
            .I(N__2342));
    InMux I__262 (
            .O(N__2345),
            .I(N__2339));
    LocalMux I__261 (
            .O(N__2342),
            .I(\pulse_counter.internal_count_10 ));
    LocalMux I__260 (
            .O(N__2339),
            .I(\pulse_counter.internal_count_10 ));
    InMux I__259 (
            .O(N__2334),
            .I(\pulse_counter.n721 ));
    InMux I__258 (
            .O(N__2331),
            .I(N__2327));
    InMux I__257 (
            .O(N__2330),
            .I(N__2324));
    LocalMux I__256 (
            .O(N__2327),
            .I(\pulse_counter.internal_count_11 ));
    LocalMux I__255 (
            .O(N__2324),
            .I(\pulse_counter.internal_count_11 ));
    InMux I__254 (
            .O(N__2319),
            .I(\pulse_counter.n722 ));
    InMux I__253 (
            .O(N__2316),
            .I(N__2312));
    InMux I__252 (
            .O(N__2315),
            .I(N__2309));
    LocalMux I__251 (
            .O(N__2312),
            .I(\pulse_counter.internal_count_12 ));
    LocalMux I__250 (
            .O(N__2309),
            .I(\pulse_counter.internal_count_12 ));
    InMux I__249 (
            .O(N__2304),
            .I(\pulse_counter.n723 ));
    InMux I__248 (
            .O(N__2301),
            .I(N__2297));
    InMux I__247 (
            .O(N__2300),
            .I(N__2294));
    LocalMux I__246 (
            .O(N__2297),
            .I(\pulse_counter.internal_count_13 ));
    LocalMux I__245 (
            .O(N__2294),
            .I(\pulse_counter.internal_count_13 ));
    InMux I__244 (
            .O(N__2289),
            .I(\pulse_counter.n724 ));
    CascadeMux I__243 (
            .O(N__2286),
            .I(N__2283));
    InMux I__242 (
            .O(N__2283),
            .I(N__2277));
    InMux I__241 (
            .O(N__2282),
            .I(N__2277));
    LocalMux I__240 (
            .O(N__2277),
            .I(N__2274));
    Span12Mux_h I__239 (
            .O(N__2274),
            .I(N__2271));
    Span12Mux_v I__238 (
            .O(N__2271),
            .I(N__2268));
    Odrv12 I__237 (
            .O(N__2268),
            .I(divide_enable_c));
    CEMux I__236 (
            .O(N__2265),
            .I(N__2262));
    LocalMux I__235 (
            .O(N__2262),
            .I(N__2258));
    CEMux I__234 (
            .O(N__2261),
            .I(N__2255));
    Span4Mux_v I__233 (
            .O(N__2258),
            .I(N__2250));
    LocalMux I__232 (
            .O(N__2255),
            .I(N__2250));
    Span4Mux_h I__231 (
            .O(N__2250),
            .I(N__2247));
    Odrv4 I__230 (
            .O(N__2247),
            .I(n176));
    InMux I__229 (
            .O(N__2244),
            .I(N__2240));
    InMux I__228 (
            .O(N__2243),
            .I(N__2237));
    LocalMux I__227 (
            .O(N__2240),
            .I(output_state));
    LocalMux I__226 (
            .O(N__2237),
            .I(output_state));
    InMux I__225 (
            .O(N__2232),
            .I(N__2229));
    LocalMux I__224 (
            .O(N__2229),
            .I(N__2226));
    Span4Mux_v I__223 (
            .O(N__2226),
            .I(N__2223));
    Span4Mux_v I__222 (
            .O(N__2223),
            .I(N__2220));
    Sp12to4 I__221 (
            .O(N__2220),
            .I(N__2217));
    Odrv12 I__220 (
            .O(N__2217),
            .I(constant_v_c));
    InMux I__219 (
            .O(N__2214),
            .I(N__2210));
    InMux I__218 (
            .O(N__2213),
            .I(N__2207));
    LocalMux I__217 (
            .O(N__2210),
            .I(\pulse_counter.internal_count_0 ));
    LocalMux I__216 (
            .O(N__2207),
            .I(\pulse_counter.internal_count_0 ));
    InMux I__215 (
            .O(N__2202),
            .I(bfn_2_7_0_));
    InMux I__214 (
            .O(N__2199),
            .I(N__2195));
    InMux I__213 (
            .O(N__2198),
            .I(N__2192));
    LocalMux I__212 (
            .O(N__2195),
            .I(\pulse_counter.internal_count_1 ));
    LocalMux I__211 (
            .O(N__2192),
            .I(\pulse_counter.internal_count_1 ));
    InMux I__210 (
            .O(N__2187),
            .I(\pulse_counter.n712 ));
    InMux I__209 (
            .O(N__2184),
            .I(N__2180));
    InMux I__208 (
            .O(N__2183),
            .I(N__2177));
    LocalMux I__207 (
            .O(N__2180),
            .I(\pulse_counter.internal_count_2 ));
    LocalMux I__206 (
            .O(N__2177),
            .I(\pulse_counter.internal_count_2 ));
    InMux I__205 (
            .O(N__2172),
            .I(\pulse_counter.n713 ));
    InMux I__204 (
            .O(N__2169),
            .I(N__2165));
    InMux I__203 (
            .O(N__2168),
            .I(N__2162));
    LocalMux I__202 (
            .O(N__2165),
            .I(\pulse_counter.internal_count_3 ));
    LocalMux I__201 (
            .O(N__2162),
            .I(\pulse_counter.internal_count_3 ));
    InMux I__200 (
            .O(N__2157),
            .I(\pulse_counter.n714 ));
    InMux I__199 (
            .O(N__2154),
            .I(N__2150));
    InMux I__198 (
            .O(N__2153),
            .I(N__2147));
    LocalMux I__197 (
            .O(N__2150),
            .I(\pulse_counter.internal_count_4 ));
    LocalMux I__196 (
            .O(N__2147),
            .I(\pulse_counter.internal_count_4 ));
    InMux I__195 (
            .O(N__2142),
            .I(\pulse_counter.n715 ));
    InMux I__194 (
            .O(N__2139),
            .I(\pulse_counter.n734 ));
    InMux I__193 (
            .O(N__2136),
            .I(bfn_1_8_0_));
    InMux I__192 (
            .O(N__2133),
            .I(\pulse_counter.n736 ));
    InMux I__191 (
            .O(N__2130),
            .I(\pulse_counter.n737 ));
    InMux I__190 (
            .O(N__2127),
            .I(\pulse_counter.n738 ));
    InMux I__189 (
            .O(N__2124),
            .I(\pulse_counter.n739 ));
    InMux I__188 (
            .O(N__2121),
            .I(\pulse_counter.n740 ));
    InMux I__187 (
            .O(N__2118),
            .I(\pulse_counter.n741 ));
    InMux I__186 (
            .O(N__2115),
            .I(\pulse_counter.n742 ));
    InMux I__185 (
            .O(N__2112),
            .I(bfn_1_7_0_));
    InMux I__184 (
            .O(N__2109),
            .I(\pulse_counter.n728 ));
    InMux I__183 (
            .O(N__2106),
            .I(\pulse_counter.n729 ));
    InMux I__182 (
            .O(N__2103),
            .I(\pulse_counter.n730 ));
    InMux I__181 (
            .O(N__2100),
            .I(\pulse_counter.n731 ));
    InMux I__180 (
            .O(N__2097),
            .I(\pulse_counter.n732 ));
    InMux I__179 (
            .O(N__2094),
            .I(\pulse_counter.n733 ));
    defparam IN_MUX_bfv_6_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_7_0_));
    defparam IN_MUX_bfv_6_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_8_0_ (
            .carryinitin(\row_counter.n703 ),
            .carryinitout(bfn_6_8_0_));
    defparam IN_MUX_bfv_6_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_9_0_ (
            .carryinitin(\row_counter.n711 ),
            .carryinitout(bfn_6_9_0_));
    defparam IN_MUX_bfv_5_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_7_0_));
    defparam IN_MUX_bfv_5_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_8_0_ (
            .carryinitin(\row_counter.n750 ),
            .carryinitout(bfn_5_8_0_));
    defparam IN_MUX_bfv_2_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_7_0_));
    defparam IN_MUX_bfv_2_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_8_0_ (
            .carryinitin(\pulse_counter.n719 ),
            .carryinitout(bfn_2_8_0_));
    defparam IN_MUX_bfv_2_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_9_0_ (
            .carryinitin(\pulse_counter.n727 ),
            .carryinitout(bfn_2_9_0_));
    defparam IN_MUX_bfv_1_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_7_0_));
    defparam IN_MUX_bfv_1_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_8_0_ (
            .carryinitin(\pulse_counter.n735 ),
            .carryinitout(bfn_1_8_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \pulse_counter.internal_count__i0_LC_1_7_0 .C_ON=1'b1;
    defparam \pulse_counter.internal_count__i0_LC_1_7_0 .SEQ_MODE=4'b1000;
    defparam \pulse_counter.internal_count__i0_LC_1_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pulse_counter.internal_count__i0_LC_1_7_0  (
            .in0(_gnd_net_),
            .in1(N__2213),
            .in2(_gnd_net_),
            .in3(N__2112),
            .lcout(\pulse_counter.internal_count_0 ),
            .ltout(),
            .carryin(bfn_1_7_0_),
            .carryout(\pulse_counter.n728 ),
            .clk(N__2631),
            .ce(N__2265),
            .sr(N__3919));
    defparam \pulse_counter.internal_count__i1_LC_1_7_1 .C_ON=1'b1;
    defparam \pulse_counter.internal_count__i1_LC_1_7_1 .SEQ_MODE=4'b1000;
    defparam \pulse_counter.internal_count__i1_LC_1_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pulse_counter.internal_count__i1_LC_1_7_1  (
            .in0(_gnd_net_),
            .in1(N__2198),
            .in2(_gnd_net_),
            .in3(N__2109),
            .lcout(\pulse_counter.internal_count_1 ),
            .ltout(),
            .carryin(\pulse_counter.n728 ),
            .carryout(\pulse_counter.n729 ),
            .clk(N__2631),
            .ce(N__2265),
            .sr(N__3919));
    defparam \pulse_counter.internal_count__i2_LC_1_7_2 .C_ON=1'b1;
    defparam \pulse_counter.internal_count__i2_LC_1_7_2 .SEQ_MODE=4'b1000;
    defparam \pulse_counter.internal_count__i2_LC_1_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pulse_counter.internal_count__i2_LC_1_7_2  (
            .in0(_gnd_net_),
            .in1(N__2184),
            .in2(_gnd_net_),
            .in3(N__2106),
            .lcout(\pulse_counter.internal_count_2 ),
            .ltout(),
            .carryin(\pulse_counter.n729 ),
            .carryout(\pulse_counter.n730 ),
            .clk(N__2631),
            .ce(N__2265),
            .sr(N__3919));
    defparam \pulse_counter.internal_count__i3_LC_1_7_3 .C_ON=1'b1;
    defparam \pulse_counter.internal_count__i3_LC_1_7_3 .SEQ_MODE=4'b1000;
    defparam \pulse_counter.internal_count__i3_LC_1_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pulse_counter.internal_count__i3_LC_1_7_3  (
            .in0(_gnd_net_),
            .in1(N__2169),
            .in2(_gnd_net_),
            .in3(N__2103),
            .lcout(\pulse_counter.internal_count_3 ),
            .ltout(),
            .carryin(\pulse_counter.n730 ),
            .carryout(\pulse_counter.n731 ),
            .clk(N__2631),
            .ce(N__2265),
            .sr(N__3919));
    defparam \pulse_counter.internal_count__i4_LC_1_7_4 .C_ON=1'b1;
    defparam \pulse_counter.internal_count__i4_LC_1_7_4 .SEQ_MODE=4'b1000;
    defparam \pulse_counter.internal_count__i4_LC_1_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pulse_counter.internal_count__i4_LC_1_7_4  (
            .in0(_gnd_net_),
            .in1(N__2154),
            .in2(_gnd_net_),
            .in3(N__2100),
            .lcout(\pulse_counter.internal_count_4 ),
            .ltout(),
            .carryin(\pulse_counter.n731 ),
            .carryout(\pulse_counter.n732 ),
            .clk(N__2631),
            .ce(N__2265),
            .sr(N__3919));
    defparam \pulse_counter.internal_count__i5_LC_1_7_5 .C_ON=1'b1;
    defparam \pulse_counter.internal_count__i5_LC_1_7_5 .SEQ_MODE=4'b1000;
    defparam \pulse_counter.internal_count__i5_LC_1_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pulse_counter.internal_count__i5_LC_1_7_5  (
            .in0(_gnd_net_),
            .in1(N__2421),
            .in2(_gnd_net_),
            .in3(N__2097),
            .lcout(\pulse_counter.internal_count_5 ),
            .ltout(),
            .carryin(\pulse_counter.n732 ),
            .carryout(\pulse_counter.n733 ),
            .clk(N__2631),
            .ce(N__2265),
            .sr(N__3919));
    defparam \pulse_counter.internal_count__i6_LC_1_7_6 .C_ON=1'b1;
    defparam \pulse_counter.internal_count__i6_LC_1_7_6 .SEQ_MODE=4'b1000;
    defparam \pulse_counter.internal_count__i6_LC_1_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pulse_counter.internal_count__i6_LC_1_7_6  (
            .in0(_gnd_net_),
            .in1(N__2406),
            .in2(_gnd_net_),
            .in3(N__2094),
            .lcout(\pulse_counter.internal_count_6 ),
            .ltout(),
            .carryin(\pulse_counter.n733 ),
            .carryout(\pulse_counter.n734 ),
            .clk(N__2631),
            .ce(N__2265),
            .sr(N__3919));
    defparam \pulse_counter.internal_count__i7_LC_1_7_7 .C_ON=1'b1;
    defparam \pulse_counter.internal_count__i7_LC_1_7_7 .SEQ_MODE=4'b1000;
    defparam \pulse_counter.internal_count__i7_LC_1_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pulse_counter.internal_count__i7_LC_1_7_7  (
            .in0(_gnd_net_),
            .in1(N__2391),
            .in2(_gnd_net_),
            .in3(N__2139),
            .lcout(\pulse_counter.internal_count_7 ),
            .ltout(),
            .carryin(\pulse_counter.n734 ),
            .carryout(\pulse_counter.n735 ),
            .clk(N__2631),
            .ce(N__2265),
            .sr(N__3919));
    defparam \pulse_counter.internal_count__i8_LC_1_8_0 .C_ON=1'b1;
    defparam \pulse_counter.internal_count__i8_LC_1_8_0 .SEQ_MODE=4'b1000;
    defparam \pulse_counter.internal_count__i8_LC_1_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pulse_counter.internal_count__i8_LC_1_8_0  (
            .in0(_gnd_net_),
            .in1(N__2376),
            .in2(_gnd_net_),
            .in3(N__2136),
            .lcout(\pulse_counter.internal_count_8 ),
            .ltout(),
            .carryin(bfn_1_8_0_),
            .carryout(\pulse_counter.n736 ),
            .clk(N__2629),
            .ce(N__2261),
            .sr(N__3915));
    defparam \pulse_counter.internal_count__i9_LC_1_8_1 .C_ON=1'b1;
    defparam \pulse_counter.internal_count__i9_LC_1_8_1 .SEQ_MODE=4'b1000;
    defparam \pulse_counter.internal_count__i9_LC_1_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pulse_counter.internal_count__i9_LC_1_8_1  (
            .in0(_gnd_net_),
            .in1(N__2361),
            .in2(_gnd_net_),
            .in3(N__2133),
            .lcout(\pulse_counter.internal_count_9 ),
            .ltout(),
            .carryin(\pulse_counter.n736 ),
            .carryout(\pulse_counter.n737 ),
            .clk(N__2629),
            .ce(N__2261),
            .sr(N__3915));
    defparam \pulse_counter.internal_count__i10_LC_1_8_2 .C_ON=1'b1;
    defparam \pulse_counter.internal_count__i10_LC_1_8_2 .SEQ_MODE=4'b1000;
    defparam \pulse_counter.internal_count__i10_LC_1_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pulse_counter.internal_count__i10_LC_1_8_2  (
            .in0(_gnd_net_),
            .in1(N__2346),
            .in2(_gnd_net_),
            .in3(N__2130),
            .lcout(\pulse_counter.internal_count_10 ),
            .ltout(),
            .carryin(\pulse_counter.n737 ),
            .carryout(\pulse_counter.n738 ),
            .clk(N__2629),
            .ce(N__2261),
            .sr(N__3915));
    defparam \pulse_counter.internal_count__i11_LC_1_8_3 .C_ON=1'b1;
    defparam \pulse_counter.internal_count__i11_LC_1_8_3 .SEQ_MODE=4'b1000;
    defparam \pulse_counter.internal_count__i11_LC_1_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pulse_counter.internal_count__i11_LC_1_8_3  (
            .in0(_gnd_net_),
            .in1(N__2331),
            .in2(_gnd_net_),
            .in3(N__2127),
            .lcout(\pulse_counter.internal_count_11 ),
            .ltout(),
            .carryin(\pulse_counter.n738 ),
            .carryout(\pulse_counter.n739 ),
            .clk(N__2629),
            .ce(N__2261),
            .sr(N__3915));
    defparam \pulse_counter.internal_count__i12_LC_1_8_4 .C_ON=1'b1;
    defparam \pulse_counter.internal_count__i12_LC_1_8_4 .SEQ_MODE=4'b1000;
    defparam \pulse_counter.internal_count__i12_LC_1_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pulse_counter.internal_count__i12_LC_1_8_4  (
            .in0(_gnd_net_),
            .in1(N__2316),
            .in2(_gnd_net_),
            .in3(N__2124),
            .lcout(\pulse_counter.internal_count_12 ),
            .ltout(),
            .carryin(\pulse_counter.n739 ),
            .carryout(\pulse_counter.n740 ),
            .clk(N__2629),
            .ce(N__2261),
            .sr(N__3915));
    defparam \pulse_counter.internal_count__i13_LC_1_8_5 .C_ON=1'b1;
    defparam \pulse_counter.internal_count__i13_LC_1_8_5 .SEQ_MODE=4'b1000;
    defparam \pulse_counter.internal_count__i13_LC_1_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pulse_counter.internal_count__i13_LC_1_8_5  (
            .in0(_gnd_net_),
            .in1(N__2301),
            .in2(_gnd_net_),
            .in3(N__2121),
            .lcout(\pulse_counter.internal_count_13 ),
            .ltout(),
            .carryin(\pulse_counter.n740 ),
            .carryout(\pulse_counter.n741 ),
            .clk(N__2629),
            .ce(N__2261),
            .sr(N__3915));
    defparam \pulse_counter.internal_count__i14_LC_1_8_6 .C_ON=1'b1;
    defparam \pulse_counter.internal_count__i14_LC_1_8_6 .SEQ_MODE=4'b1000;
    defparam \pulse_counter.internal_count__i14_LC_1_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pulse_counter.internal_count__i14_LC_1_8_6  (
            .in0(_gnd_net_),
            .in1(N__2540),
            .in2(_gnd_net_),
            .in3(N__2118),
            .lcout(\pulse_counter.internal_count_14 ),
            .ltout(),
            .carryin(\pulse_counter.n741 ),
            .carryout(\pulse_counter.n742 ),
            .clk(N__2629),
            .ce(N__2261),
            .sr(N__3915));
    defparam \pulse_counter.internal_count__i15_LC_1_8_7 .C_ON=1'b0;
    defparam \pulse_counter.internal_count__i15_LC_1_8_7 .SEQ_MODE=4'b1000;
    defparam \pulse_counter.internal_count__i15_LC_1_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pulse_counter.internal_count__i15_LC_1_8_7  (
            .in0(_gnd_net_),
            .in1(N__2522),
            .in2(_gnd_net_),
            .in3(N__2115),
            .lcout(\pulse_counter.internal_count_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2629),
            .ce(N__2261),
            .sr(N__3915));
    defparam output_state_20_LC_1_9_2.C_ON=1'b0;
    defparam output_state_20_LC_1_9_2.SEQ_MODE=4'b1000;
    defparam output_state_20_LC_1_9_2.LUT_INIT=16'b1010101001100010;
    LogicCell40 output_state_20_LC_1_9_2 (
            .in0(N__2243),
            .in1(N__2647),
            .in2(N__2286),
            .in3(N__3878),
            .lcout(output_state),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2628),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_LC_1_9_6.C_ON=1'b0;
    defparam i1_3_lut_LC_1_9_6.SEQ_MODE=4'b0000;
    defparam i1_3_lut_LC_1_9_6.LUT_INIT=16'b1111111100100010;
    LogicCell40 i1_3_lut_LC_1_9_6 (
            .in0(N__2282),
            .in1(N__2646),
            .in2(_gnd_net_),
            .in3(N__3877),
            .lcout(n176),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam output_state_I_0_21_2_lut_LC_1_10_6.C_ON=1'b0;
    defparam output_state_I_0_21_2_lut_LC_1_10_6.SEQ_MODE=4'b0000;
    defparam output_state_I_0_21_2_lut_LC_1_10_6.LUT_INIT=16'b1010101000000000;
    LogicCell40 output_state_I_0_21_2_lut_LC_1_10_6 (
            .in0(N__2244),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2232),
            .lcout(divided_pulse_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pulse_counter.sub_8_add_2_2_lut_LC_2_7_0 .C_ON=1'b1;
    defparam \pulse_counter.sub_8_add_2_2_lut_LC_2_7_0 .SEQ_MODE=4'b0000;
    defparam \pulse_counter.sub_8_add_2_2_lut_LC_2_7_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pulse_counter.sub_8_add_2_2_lut_LC_2_7_0  (
            .in0(N__2214),
            .in1(N__2577),
            .in2(_gnd_net_),
            .in3(N__2202),
            .lcout(n1_adj_117),
            .ltout(),
            .carryin(bfn_2_7_0_),
            .carryout(\pulse_counter.n712 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pulse_counter.sub_8_add_2_3_lut_LC_2_7_1 .C_ON=1'b1;
    defparam \pulse_counter.sub_8_add_2_3_lut_LC_2_7_1 .SEQ_MODE=4'b0000;
    defparam \pulse_counter.sub_8_add_2_3_lut_LC_2_7_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pulse_counter.sub_8_add_2_3_lut_LC_2_7_1  (
            .in0(N__2199),
            .in1(N__2550),
            .in2(N__4218),
            .in3(N__2187),
            .lcout(n2_adj_99),
            .ltout(),
            .carryin(\pulse_counter.n712 ),
            .carryout(\pulse_counter.n713 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pulse_counter.sub_8_add_2_4_lut_LC_2_7_2 .C_ON=1'b1;
    defparam \pulse_counter.sub_8_add_2_4_lut_LC_2_7_2 .SEQ_MODE=4'b0000;
    defparam \pulse_counter.sub_8_add_2_4_lut_LC_2_7_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pulse_counter.sub_8_add_2_4_lut_LC_2_7_2  (
            .in0(N__2183),
            .in1(N__4201),
            .in2(N__2613),
            .in3(N__2172),
            .lcout(n3_adj_118),
            .ltout(),
            .carryin(\pulse_counter.n713 ),
            .carryout(\pulse_counter.n714 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pulse_counter.sub_8_add_2_5_lut_LC_2_7_3 .C_ON=1'b1;
    defparam \pulse_counter.sub_8_add_2_5_lut_LC_2_7_3 .SEQ_MODE=4'b0000;
    defparam \pulse_counter.sub_8_add_2_5_lut_LC_2_7_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pulse_counter.sub_8_add_2_5_lut_LC_2_7_3  (
            .in0(N__2168),
            .in1(N__2568),
            .in2(N__4219),
            .in3(N__2157),
            .lcout(n4_adj_116),
            .ltout(),
            .carryin(\pulse_counter.n714 ),
            .carryout(\pulse_counter.n715 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pulse_counter.sub_8_add_2_6_lut_LC_2_7_4 .C_ON=1'b1;
    defparam \pulse_counter.sub_8_add_2_6_lut_LC_2_7_4 .SEQ_MODE=4'b0000;
    defparam \pulse_counter.sub_8_add_2_6_lut_LC_2_7_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pulse_counter.sub_8_add_2_6_lut_LC_2_7_4  (
            .in0(N__2153),
            .in1(N__4205),
            .in2(N__2739),
            .in3(N__2142),
            .lcout(n5_adj_120),
            .ltout(),
            .carryin(\pulse_counter.n715 ),
            .carryout(\pulse_counter.n716 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pulse_counter.sub_8_add_2_7_lut_LC_2_7_5 .C_ON=1'b1;
    defparam \pulse_counter.sub_8_add_2_7_lut_LC_2_7_5 .SEQ_MODE=4'b0000;
    defparam \pulse_counter.sub_8_add_2_7_lut_LC_2_7_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pulse_counter.sub_8_add_2_7_lut_LC_2_7_5  (
            .in0(N__2420),
            .in1(N__2727),
            .in2(N__4220),
            .in3(N__2409),
            .lcout(n6_adj_119),
            .ltout(),
            .carryin(\pulse_counter.n716 ),
            .carryout(\pulse_counter.n717 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pulse_counter.sub_8_add_2_8_lut_LC_2_7_6 .C_ON=1'b1;
    defparam \pulse_counter.sub_8_add_2_8_lut_LC_2_7_6 .SEQ_MODE=4'b0000;
    defparam \pulse_counter.sub_8_add_2_8_lut_LC_2_7_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pulse_counter.sub_8_add_2_8_lut_LC_2_7_6  (
            .in0(N__2405),
            .in1(N__2757),
            .in2(N__4212),
            .in3(N__2394),
            .lcout(n7),
            .ltout(),
            .carryin(\pulse_counter.n717 ),
            .carryout(\pulse_counter.n718 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pulse_counter.sub_8_add_2_9_lut_LC_2_7_7 .C_ON=1'b1;
    defparam \pulse_counter.sub_8_add_2_9_lut_LC_2_7_7 .SEQ_MODE=4'b0000;
    defparam \pulse_counter.sub_8_add_2_9_lut_LC_2_7_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pulse_counter.sub_8_add_2_9_lut_LC_2_7_7  (
            .in0(N__2390),
            .in1(N__2706),
            .in2(N__4221),
            .in3(N__2379),
            .lcout(n8),
            .ltout(),
            .carryin(\pulse_counter.n718 ),
            .carryout(\pulse_counter.n719 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pulse_counter.sub_8_add_2_10_lut_LC_2_8_0 .C_ON=1'b1;
    defparam \pulse_counter.sub_8_add_2_10_lut_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \pulse_counter.sub_8_add_2_10_lut_LC_2_8_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pulse_counter.sub_8_add_2_10_lut_LC_2_8_0  (
            .in0(N__2375),
            .in1(N__2718),
            .in2(N__4213),
            .in3(N__2364),
            .lcout(n9),
            .ltout(),
            .carryin(bfn_2_8_0_),
            .carryout(\pulse_counter.n720 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pulse_counter.sub_8_add_2_11_lut_LC_2_8_1 .C_ON=1'b1;
    defparam \pulse_counter.sub_8_add_2_11_lut_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \pulse_counter.sub_8_add_2_11_lut_LC_2_8_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pulse_counter.sub_8_add_2_11_lut_LC_2_8_1  (
            .in0(N__2360),
            .in1(N__2748),
            .in2(N__4216),
            .in3(N__2349),
            .lcout(n10),
            .ltout(),
            .carryin(\pulse_counter.n720 ),
            .carryout(\pulse_counter.n721 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pulse_counter.sub_8_add_2_12_lut_LC_2_8_2 .C_ON=1'b1;
    defparam \pulse_counter.sub_8_add_2_12_lut_LC_2_8_2 .SEQ_MODE=4'b0000;
    defparam \pulse_counter.sub_8_add_2_12_lut_LC_2_8_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pulse_counter.sub_8_add_2_12_lut_LC_2_8_2  (
            .in0(N__2345),
            .in1(N__2766),
            .in2(N__4214),
            .in3(N__2334),
            .lcout(n11),
            .ltout(),
            .carryin(\pulse_counter.n721 ),
            .carryout(\pulse_counter.n722 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pulse_counter.sub_8_add_2_13_lut_LC_2_8_3 .C_ON=1'b1;
    defparam \pulse_counter.sub_8_add_2_13_lut_LC_2_8_3 .SEQ_MODE=4'b0000;
    defparam \pulse_counter.sub_8_add_2_13_lut_LC_2_8_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pulse_counter.sub_8_add_2_13_lut_LC_2_8_3  (
            .in0(N__2330),
            .in1(N__2427),
            .in2(N__4217),
            .in3(N__2319),
            .lcout(n12),
            .ltout(),
            .carryin(\pulse_counter.n722 ),
            .carryout(\pulse_counter.n723 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pulse_counter.sub_8_add_2_14_lut_LC_2_8_4 .C_ON=1'b1;
    defparam \pulse_counter.sub_8_add_2_14_lut_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \pulse_counter.sub_8_add_2_14_lut_LC_2_8_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pulse_counter.sub_8_add_2_14_lut_LC_2_8_4  (
            .in0(N__2315),
            .in1(N__2559),
            .in2(N__4215),
            .in3(N__2304),
            .lcout(\pulse_counter.n13 ),
            .ltout(),
            .carryin(\pulse_counter.n723 ),
            .carryout(\pulse_counter.n724 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pulse_counter.sub_8_add_2_15_lut_LC_2_8_5 .C_ON=1'b1;
    defparam \pulse_counter.sub_8_add_2_15_lut_LC_2_8_5 .SEQ_MODE=4'b0000;
    defparam \pulse_counter.sub_8_add_2_15_lut_LC_2_8_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pulse_counter.sub_8_add_2_15_lut_LC_2_8_5  (
            .in0(N__2300),
            .in1(N__4189),
            .in2(N__2658),
            .in3(N__2289),
            .lcout(n14),
            .ltout(),
            .carryin(\pulse_counter.n724 ),
            .carryout(\pulse_counter.n725 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pulse_counter.sub_8_add_2_16_lut_LC_2_8_6 .C_ON=1'b1;
    defparam \pulse_counter.sub_8_add_2_16_lut_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \pulse_counter.sub_8_add_2_16_lut_LC_2_8_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pulse_counter.sub_8_add_2_16_lut_LC_2_8_6  (
            .in0(N__2541),
            .in1(N__4197),
            .in2(N__2601),
            .in3(N__2526),
            .lcout(n15),
            .ltout(),
            .carryin(\pulse_counter.n725 ),
            .carryout(\pulse_counter.n726 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pulse_counter.sub_8_add_2_17_lut_LC_2_8_7 .C_ON=1'b1;
    defparam \pulse_counter.sub_8_add_2_17_lut_LC_2_8_7 .SEQ_MODE=4'b0000;
    defparam \pulse_counter.sub_8_add_2_17_lut_LC_2_8_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pulse_counter.sub_8_add_2_17_lut_LC_2_8_7  (
            .in0(N__2523),
            .in1(N__4190),
            .in2(N__2589),
            .in3(N__2508),
            .lcout(n16),
            .ltout(),
            .carryin(\pulse_counter.n726 ),
            .carryout(\pulse_counter.n727 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pulse_counter.sub_8_add_2_18_lut_LC_2_9_0 .C_ON=1'b0;
    defparam \pulse_counter.sub_8_add_2_18_lut_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \pulse_counter.sub_8_add_2_18_lut_LC_2_9_0 .LUT_INIT=16'b1110110111011110;
    LogicCell40 \pulse_counter.sub_8_add_2_18_lut_LC_2_9_0  (
            .in0(N__4119),
            .in1(N__2505),
            .in2(_gnd_net_),
            .in3(N__2499),
            .lcout(n787),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i732_2_lut_LC_2_9_1.C_ON=1'b0;
    defparam i732_2_lut_LC_2_9_1.SEQ_MODE=4'b0000;
    defparam i732_2_lut_LC_2_9_1.LUT_INIT=16'b1111111111001100;
    LogicCell40 i732_2_lut_LC_2_9_1 (
            .in0(_gnd_net_),
            .in1(N__2496),
            .in2(_gnd_net_),
            .in3(N__2487),
            .lcout(),
            .ltout(n795_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i754_4_lut_LC_2_9_2.C_ON=1'b0;
    defparam i754_4_lut_LC_2_9_2.SEQ_MODE=4'b0000;
    defparam i754_4_lut_LC_2_9_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i754_4_lut_LC_2_9_2 (
            .in0(N__2478),
            .in1(N__2469),
            .in2(N__2463),
            .in3(N__2460),
            .lcout(),
            .ltout(n817_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i762_4_lut_LC_2_9_3.C_ON=1'b0;
    defparam i762_4_lut_LC_2_9_3.SEQ_MODE=4'b0000;
    defparam i762_4_lut_LC_2_9_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i762_4_lut_LC_2_9_3 (
            .in0(N__2451),
            .in1(N__2445),
            .in2(N__2439),
            .in3(N__2436),
            .lcout(),
            .ltout(n825_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pulse_counter.internal_count_reached_18_LC_2_9_4 .C_ON=1'b0;
    defparam \pulse_counter.internal_count_reached_18_LC_2_9_4 .SEQ_MODE=4'b1000;
    defparam \pulse_counter.internal_count_reached_18_LC_2_9_4 .LUT_INIT=16'b0000000010101011;
    LogicCell40 \pulse_counter.internal_count_reached_18_LC_2_9_4  (
            .in0(N__2649),
            .in1(N__2883),
            .in2(N__2430),
            .in3(N__3879),
            .lcout(count_done),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2630),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.output_enable_I_0_i12_2_lut_LC_2_9_5 .C_ON=1'b0;
    defparam \divider_sr.output_enable_I_0_i12_2_lut_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \divider_sr.output_enable_I_0_i12_2_lut_LC_2_9_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \divider_sr.output_enable_I_0_i12_2_lut_LC_2_9_5  (
            .in0(N__2781),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4622),
            .lcout(sr_divider_data_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.output_enable_I_0_i14_2_lut_LC_2_9_6 .C_ON=1'b0;
    defparam \divider_sr.output_enable_I_0_i14_2_lut_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \divider_sr.output_enable_I_0_i14_2_lut_LC_2_9_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \divider_sr.output_enable_I_0_i14_2_lut_LC_2_9_6  (
            .in0(N__4623),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3027),
            .lcout(sr_divider_data_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam reset_signal_19_LC_2_9_7.C_ON=1'b0;
    defparam reset_signal_19_LC_2_9_7.SEQ_MODE=4'b1000;
    defparam reset_signal_19_LC_2_9_7.LUT_INIT=16'b1111111101000100;
    LogicCell40 reset_signal_19_LC_2_9_7 (
            .in0(N__3880),
            .in1(N__2648),
            .in2(_gnd_net_),
            .in3(N__3828),
            .lcout(reset_signal),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2630),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.output_enable_I_0_i3_2_lut_LC_2_10_0 .C_ON=1'b0;
    defparam \divider_sr.output_enable_I_0_i3_2_lut_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \divider_sr.output_enable_I_0_i3_2_lut_LC_2_10_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \divider_sr.output_enable_I_0_i3_2_lut_LC_2_10_0  (
            .in0(N__4591),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3350),
            .lcout(sr_divider_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.output_enable_I_0_i15_2_lut_LC_2_10_1 .C_ON=1'b0;
    defparam \divider_sr.output_enable_I_0_i15_2_lut_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \divider_sr.output_enable_I_0_i15_2_lut_LC_2_10_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \divider_sr.output_enable_I_0_i15_2_lut_LC_2_10_1  (
            .in0(_gnd_net_),
            .in1(N__4587),
            .in2(_gnd_net_),
            .in3(N__2808),
            .lcout(sr_divider_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.output_enable_I_0_i16_2_lut_LC_2_10_2 .C_ON=1'b0;
    defparam \divider_sr.output_enable_I_0_i16_2_lut_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \divider_sr.output_enable_I_0_i16_2_lut_LC_2_10_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \divider_sr.output_enable_I_0_i16_2_lut_LC_2_10_2  (
            .in0(N__4588),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2793),
            .lcout(sr_divider_data_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.output_enable_I_0_i1_2_lut_LC_2_10_3 .C_ON=1'b0;
    defparam \divider_sr.output_enable_I_0_i1_2_lut_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \divider_sr.output_enable_I_0_i1_2_lut_LC_2_10_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \divider_sr.output_enable_I_0_i1_2_lut_LC_2_10_3  (
            .in0(_gnd_net_),
            .in1(N__4589),
            .in2(_gnd_net_),
            .in3(N__3393),
            .lcout(sr_divider_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.output_enable_I_0_i4_2_lut_LC_2_10_4 .C_ON=1'b0;
    defparam \divider_sr.output_enable_I_0_i4_2_lut_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \divider_sr.output_enable_I_0_i4_2_lut_LC_2_10_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \divider_sr.output_enable_I_0_i4_2_lut_LC_2_10_4  (
            .in0(N__4592),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3165),
            .lcout(sr_divider_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.output_enable_I_0_i13_2_lut_LC_2_10_5 .C_ON=1'b0;
    defparam \divider_sr.output_enable_I_0_i13_2_lut_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \divider_sr.output_enable_I_0_i13_2_lut_LC_2_10_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \divider_sr.output_enable_I_0_i13_2_lut_LC_2_10_5  (
            .in0(N__3047),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4586),
            .lcout(sr_divider_data_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.output_enable_I_0_i2_2_lut_LC_2_10_6 .C_ON=1'b0;
    defparam \divider_sr.output_enable_I_0_i2_2_lut_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \divider_sr.output_enable_I_0_i2_2_lut_LC_2_10_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \divider_sr.output_enable_I_0_i2_2_lut_LC_2_10_6  (
            .in0(N__4590),
            .in1(N__3375),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sr_divider_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.output_enable_I_0_i11_2_lut_LC_2_10_7 .C_ON=1'b0;
    defparam \divider_sr.output_enable_I_0_i11_2_lut_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \divider_sr.output_enable_I_0_i11_2_lut_LC_2_10_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \divider_sr.output_enable_I_0_i11_2_lut_LC_2_10_7  (
            .in0(_gnd_net_),
            .in1(N__4585),
            .in2(_gnd_net_),
            .in3(N__2976),
            .lcout(sr_divider_data_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.output_enable_I_0_i7_2_lut_LC_2_11_0 .C_ON=1'b0;
    defparam \divider_sr.output_enable_I_0_i7_2_lut_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \divider_sr.output_enable_I_0_i7_2_lut_LC_2_11_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \divider_sr.output_enable_I_0_i7_2_lut_LC_2_11_0  (
            .in0(N__2943),
            .in1(N__4548),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sr_divider_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.output_enable_I_0_i10_2_lut_LC_2_11_1 .C_ON=1'b0;
    defparam \divider_sr.output_enable_I_0_i10_2_lut_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \divider_sr.output_enable_I_0_i10_2_lut_LC_2_11_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \divider_sr.output_enable_I_0_i10_2_lut_LC_2_11_1  (
            .in0(N__4545),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2996),
            .lcout(sr_divider_data_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.output_enable_I_0_i5_2_lut_LC_2_11_2 .C_ON=1'b0;
    defparam \divider_sr.output_enable_I_0_i5_2_lut_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \divider_sr.output_enable_I_0_i5_2_lut_LC_2_11_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \divider_sr.output_enable_I_0_i5_2_lut_LC_2_11_2  (
            .in0(_gnd_net_),
            .in1(N__3140),
            .in2(_gnd_net_),
            .in3(N__4546),
            .lcout(sr_divider_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.output_enable_I_0_i6_2_lut_LC_2_11_4 .C_ON=1'b0;
    defparam \divider_sr.output_enable_I_0_i6_2_lut_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \divider_sr.output_enable_I_0_i6_2_lut_LC_2_11_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \divider_sr.output_enable_I_0_i6_2_lut_LC_2_11_4  (
            .in0(_gnd_net_),
            .in1(N__4547),
            .in2(_gnd_net_),
            .in3(N__2958),
            .lcout(sr_divider_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.output_enable_I_0_i9_2_lut_LC_2_11_6 .C_ON=1'b0;
    defparam \divider_sr.output_enable_I_0_i9_2_lut_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \divider_sr.output_enable_I_0_i9_2_lut_LC_2_11_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \divider_sr.output_enable_I_0_i9_2_lut_LC_2_11_6  (
            .in0(_gnd_net_),
            .in1(N__4550),
            .in2(_gnd_net_),
            .in3(N__3012),
            .lcout(sr_divider_data_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.output_enable_I_0_i8_2_lut_LC_2_11_7 .C_ON=1'b0;
    defparam \divider_sr.output_enable_I_0_i8_2_lut_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \divider_sr.output_enable_I_0_i8_2_lut_LC_2_11_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \divider_sr.output_enable_I_0_i8_2_lut_LC_2_11_7  (
            .in0(N__4549),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2927),
            .lcout(sr_divider_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i718_2_lut_LC_3_7_4.C_ON=1'b0;
    defparam i718_2_lut_LC_3_7_4.SEQ_MODE=4'b0000;
    defparam i718_2_lut_LC_3_7_4.LUT_INIT=16'b1111111111001100;
    LogicCell40 i718_2_lut_LC_3_7_4 (
            .in0(_gnd_net_),
            .in1(N__2697),
            .in2(_gnd_net_),
            .in3(N__2691),
            .lcout(n781),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i760_4_lut_LC_3_8_0.C_ON=1'b0;
    defparam i760_4_lut_LC_3_8_0.SEQ_MODE=4'b0000;
    defparam i760_4_lut_LC_3_8_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i760_4_lut_LC_3_8_0 (
            .in0(N__2685),
            .in1(N__2679),
            .in2(N__2673),
            .in3(N__2664),
            .lcout(),
            .ltout(n823_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i764_4_lut_LC_3_8_1.C_ON=1'b0;
    defparam i764_4_lut_LC_3_8_1.SEQ_MODE=4'b0000;
    defparam i764_4_lut_LC_3_8_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i764_4_lut_LC_3_8_1 (
            .in0(N__2904),
            .in1(N__2898),
            .in2(N__2892),
            .in3(N__2889),
            .lcout(n827),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i355_2_lut_3_lut_LC_3_9_2.C_ON=1'b0;
    defparam i355_2_lut_3_lut_LC_3_9_2.SEQ_MODE=4'b0000;
    defparam i355_2_lut_3_lut_LC_3_9_2.LUT_INIT=16'b0011001100100010;
    LogicCell40 i355_2_lut_3_lut_LC_3_9_2 (
            .in0(N__3892),
            .in1(N__2877),
            .in2(_gnd_net_),
            .in3(N__2836),
            .lcout(n345),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_5_LC_3_9_4.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_5_LC_3_9_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_5_LC_3_9_4.LUT_INIT=16'b1111111111101110;
    LogicCell40 i1_2_lut_3_lut_adj_5_LC_3_9_4 (
            .in0(N__3891),
            .in1(N__2876),
            .in2(_gnd_net_),
            .in3(N__2835),
            .lcout(n171),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.shifted_data_i11_LC_3_10_0 .C_ON=1'b0;
    defparam \divider_sr.shifted_data_i11_LC_3_10_0 .SEQ_MODE=4'b1000;
    defparam \divider_sr.shifted_data_i11_LC_3_10_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \divider_sr.shifted_data_i11_LC_3_10_0  (
            .in0(N__3289),
            .in1(N__2779),
            .in2(N__3236),
            .in3(N__2975),
            .lcout(shifted_data_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4708),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_LC_3_10_1.C_ON=1'b0;
    defparam i1_2_lut_3_lut_LC_3_10_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_LC_3_10_1.LUT_INIT=16'b1111111111101110;
    LogicCell40 i1_2_lut_3_lut_LC_3_10_1 (
            .in0(N__2855),
            .in1(N__2837),
            .in2(_gnd_net_),
            .in3(N__3893),
            .lcout(n169),
            .ltout(n169_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.shifted_data_i14_LC_3_10_2 .C_ON=1'b0;
    defparam \divider_sr.shifted_data_i14_LC_3_10_2 .SEQ_MODE=4'b1000;
    defparam \divider_sr.shifted_data_i14_LC_3_10_2 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \divider_sr.shifted_data_i14_LC_3_10_2  (
            .in0(N__3294),
            .in1(N__2806),
            .in2(N__2859),
            .in3(N__3026),
            .lcout(shifted_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4708),
            .ce(),
            .sr(_gnd_net_));
    defparam i340_2_lut_3_lut_LC_3_10_3.C_ON=1'b0;
    defparam i340_2_lut_3_lut_LC_3_10_3.SEQ_MODE=4'b0000;
    defparam i340_2_lut_3_lut_LC_3_10_3.LUT_INIT=16'b0101010101000100;
    LogicCell40 i340_2_lut_3_lut_LC_3_10_3 (
            .in0(N__2856),
            .in1(N__2838),
            .in2(_gnd_net_),
            .in3(N__3894),
            .lcout(n330),
            .ltout(n330_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.shifted_data_i15_LC_3_10_4 .C_ON=1'b0;
    defparam \divider_sr.shifted_data_i15_LC_3_10_4 .SEQ_MODE=4'b1000;
    defparam \divider_sr.shifted_data_i15_LC_3_10_4 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \divider_sr.shifted_data_i15_LC_3_10_4  (
            .in0(N__3211),
            .in1(N__2792),
            .in2(N__2811),
            .in3(N__2807),
            .lcout(shifted_data_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4708),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.shifted_data_i12_LC_3_10_5 .C_ON=1'b0;
    defparam \divider_sr.shifted_data_i12_LC_3_10_5 .SEQ_MODE=4'b1000;
    defparam \divider_sr.shifted_data_i12_LC_3_10_5 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \divider_sr.shifted_data_i12_LC_3_10_5  (
            .in0(N__2780),
            .in1(N__3290),
            .in2(N__3048),
            .in3(N__3210),
            .lcout(shifted_data_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4708),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.shifted_data_i13_LC_3_10_6 .C_ON=1'b0;
    defparam \divider_sr.shifted_data_i13_LC_3_10_6 .SEQ_MODE=4'b1000;
    defparam \divider_sr.shifted_data_i13_LC_3_10_6 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \divider_sr.shifted_data_i13_LC_3_10_6  (
            .in0(N__3043),
            .in1(N__3212),
            .in2(N__3315),
            .in3(N__3025),
            .lcout(shifted_data_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4708),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.shifted_data_i8_LC_3_11_0 .C_ON=1'b0;
    defparam \divider_sr.shifted_data_i8_LC_3_11_0 .SEQ_MODE=4'b1000;
    defparam \divider_sr.shifted_data_i8_LC_3_11_0 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \divider_sr.shifted_data_i8_LC_3_11_0  (
            .in0(N__2923),
            .in1(N__3221),
            .in2(N__3316),
            .in3(N__3010),
            .lcout(shifted_data_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4709),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.shifted_data_i6_LC_3_11_1 .C_ON=1'b0;
    defparam \divider_sr.shifted_data_i6_LC_3_11_1 .SEQ_MODE=4'b1000;
    defparam \divider_sr.shifted_data_i6_LC_3_11_1 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \divider_sr.shifted_data_i6_LC_3_11_1  (
            .in0(N__2956),
            .in1(N__3297),
            .in2(N__3238),
            .in3(N__2941),
            .lcout(shifted_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4709),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.shifted_data_i9_LC_3_11_2 .C_ON=1'b0;
    defparam \divider_sr.shifted_data_i9_LC_3_11_2 .SEQ_MODE=4'b1000;
    defparam \divider_sr.shifted_data_i9_LC_3_11_2 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \divider_sr.shifted_data_i9_LC_3_11_2  (
            .in0(N__3302),
            .in1(N__3222),
            .in2(N__2997),
            .in3(N__3011),
            .lcout(shifted_data_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4709),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.shifted_data_i10_LC_3_11_5 .C_ON=1'b0;
    defparam \divider_sr.shifted_data_i10_LC_3_11_5 .SEQ_MODE=4'b1000;
    defparam \divider_sr.shifted_data_i10_LC_3_11_5 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \divider_sr.shifted_data_i10_LC_3_11_5  (
            .in0(N__2992),
            .in1(N__3295),
            .in2(N__3237),
            .in3(N__2974),
            .lcout(shifted_data_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4709),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.shifted_data_i5_LC_3_11_6 .C_ON=1'b0;
    defparam \divider_sr.shifted_data_i5_LC_3_11_6 .SEQ_MODE=4'b1000;
    defparam \divider_sr.shifted_data_i5_LC_3_11_6 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \divider_sr.shifted_data_i5_LC_3_11_6  (
            .in0(N__3296),
            .in1(N__3216),
            .in2(N__3141),
            .in3(N__2957),
            .lcout(shifted_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4709),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.shifted_data_i7_LC_3_11_7 .C_ON=1'b0;
    defparam \divider_sr.shifted_data_i7_LC_3_11_7 .SEQ_MODE=4'b1000;
    defparam \divider_sr.shifted_data_i7_LC_3_11_7 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \divider_sr.shifted_data_i7_LC_3_11_7  (
            .in0(N__3220),
            .in1(N__2942),
            .in2(N__2928),
            .in3(N__3298),
            .lcout(shifted_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4709),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.shifted_data_i0_LC_5_6_3 .C_ON=1'b0;
    defparam \row_sr.shifted_data_i0_LC_5_6_3 .SEQ_MODE=4'b1000;
    defparam \row_sr.shifted_data_i0_LC_5_6_3 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \row_sr.shifted_data_i0_LC_5_6_3  (
            .in0(N__3416),
            .in1(N__4964),
            .in2(N__4878),
            .in3(N__3109),
            .lcout(shifted_data_0_adj_115),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4716),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_counter.internal_count__i0_LC_5_7_0 .C_ON=1'b1;
    defparam \row_counter.internal_count__i0_LC_5_7_0 .SEQ_MODE=4'b1000;
    defparam \row_counter.internal_count__i0_LC_5_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \row_counter.internal_count__i0_LC_5_7_0  (
            .in0(_gnd_net_),
            .in1(N__3620),
            .in2(_gnd_net_),
            .in3(N__2907),
            .lcout(\row_counter.internal_count_0 ),
            .ltout(),
            .carryin(bfn_5_7_0_),
            .carryout(\row_counter.n743 ),
            .clk(N__3803),
            .ce(N__3438),
            .sr(N__3924));
    defparam \row_counter.internal_count__i1_LC_5_7_1 .C_ON=1'b1;
    defparam \row_counter.internal_count__i1_LC_5_7_1 .SEQ_MODE=4'b1000;
    defparam \row_counter.internal_count__i1_LC_5_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \row_counter.internal_count__i1_LC_5_7_1  (
            .in0(_gnd_net_),
            .in1(N__3596),
            .in2(_gnd_net_),
            .in3(N__3075),
            .lcout(\row_counter.internal_count_1 ),
            .ltout(),
            .carryin(\row_counter.n743 ),
            .carryout(\row_counter.n744 ),
            .clk(N__3803),
            .ce(N__3438),
            .sr(N__3924));
    defparam \row_counter.internal_count__i2_LC_5_7_2 .C_ON=1'b1;
    defparam \row_counter.internal_count__i2_LC_5_7_2 .SEQ_MODE=4'b1000;
    defparam \row_counter.internal_count__i2_LC_5_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \row_counter.internal_count__i2_LC_5_7_2  (
            .in0(_gnd_net_),
            .in1(N__3573),
            .in2(_gnd_net_),
            .in3(N__3072),
            .lcout(\row_counter.internal_count_2 ),
            .ltout(),
            .carryin(\row_counter.n744 ),
            .carryout(\row_counter.n745 ),
            .clk(N__3803),
            .ce(N__3438),
            .sr(N__3924));
    defparam \row_counter.internal_count__i3_LC_5_7_3 .C_ON=1'b1;
    defparam \row_counter.internal_count__i3_LC_5_7_3 .SEQ_MODE=4'b1000;
    defparam \row_counter.internal_count__i3_LC_5_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \row_counter.internal_count__i3_LC_5_7_3  (
            .in0(_gnd_net_),
            .in1(N__3551),
            .in2(_gnd_net_),
            .in3(N__3069),
            .lcout(\row_counter.internal_count_3 ),
            .ltout(),
            .carryin(\row_counter.n745 ),
            .carryout(\row_counter.n746 ),
            .clk(N__3803),
            .ce(N__3438),
            .sr(N__3924));
    defparam \row_counter.internal_count__i4_LC_5_7_4 .C_ON=1'b1;
    defparam \row_counter.internal_count__i4_LC_5_7_4 .SEQ_MODE=4'b1000;
    defparam \row_counter.internal_count__i4_LC_5_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \row_counter.internal_count__i4_LC_5_7_4  (
            .in0(_gnd_net_),
            .in1(N__3537),
            .in2(_gnd_net_),
            .in3(N__3066),
            .lcout(\row_counter.internal_count_4 ),
            .ltout(),
            .carryin(\row_counter.n746 ),
            .carryout(\row_counter.n747 ),
            .clk(N__3803),
            .ce(N__3438),
            .sr(N__3924));
    defparam \row_counter.internal_count__i5_LC_5_7_5 .C_ON=1'b1;
    defparam \row_counter.internal_count__i5_LC_5_7_5 .SEQ_MODE=4'b1000;
    defparam \row_counter.internal_count__i5_LC_5_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \row_counter.internal_count__i5_LC_5_7_5  (
            .in0(_gnd_net_),
            .in1(N__3512),
            .in2(_gnd_net_),
            .in3(N__3063),
            .lcout(\row_counter.internal_count_5 ),
            .ltout(),
            .carryin(\row_counter.n747 ),
            .carryout(\row_counter.n748 ),
            .clk(N__3803),
            .ce(N__3438),
            .sr(N__3924));
    defparam \row_counter.internal_count__i6_LC_5_7_6 .C_ON=1'b1;
    defparam \row_counter.internal_count__i6_LC_5_7_6 .SEQ_MODE=4'b1000;
    defparam \row_counter.internal_count__i6_LC_5_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \row_counter.internal_count__i6_LC_5_7_6  (
            .in0(_gnd_net_),
            .in1(N__3498),
            .in2(_gnd_net_),
            .in3(N__3060),
            .lcout(\row_counter.internal_count_6 ),
            .ltout(),
            .carryin(\row_counter.n748 ),
            .carryout(\row_counter.n749 ),
            .clk(N__3803),
            .ce(N__3438),
            .sr(N__3924));
    defparam \row_counter.internal_count__i7_LC_5_7_7 .C_ON=1'b1;
    defparam \row_counter.internal_count__i7_LC_5_7_7 .SEQ_MODE=4'b1000;
    defparam \row_counter.internal_count__i7_LC_5_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \row_counter.internal_count__i7_LC_5_7_7  (
            .in0(_gnd_net_),
            .in1(N__3483),
            .in2(_gnd_net_),
            .in3(N__3057),
            .lcout(\row_counter.internal_count_7 ),
            .ltout(),
            .carryin(\row_counter.n749 ),
            .carryout(\row_counter.n750 ),
            .clk(N__3803),
            .ce(N__3438),
            .sr(N__3924));
    defparam \row_counter.internal_count__i8_LC_5_8_0 .C_ON=1'b1;
    defparam \row_counter.internal_count__i8_LC_5_8_0 .SEQ_MODE=4'b1000;
    defparam \row_counter.internal_count__i8_LC_5_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \row_counter.internal_count__i8_LC_5_8_0  (
            .in0(_gnd_net_),
            .in1(N__3756),
            .in2(_gnd_net_),
            .in3(N__3054),
            .lcout(\row_counter.internal_count_8 ),
            .ltout(),
            .carryin(bfn_5_8_0_),
            .carryout(\row_counter.n751 ),
            .clk(N__3802),
            .ce(N__3437),
            .sr(N__3923));
    defparam \row_counter.internal_count__i9_LC_5_8_1 .C_ON=1'b1;
    defparam \row_counter.internal_count__i9_LC_5_8_1 .SEQ_MODE=4'b1000;
    defparam \row_counter.internal_count__i9_LC_5_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \row_counter.internal_count__i9_LC_5_8_1  (
            .in0(_gnd_net_),
            .in1(N__3740),
            .in2(_gnd_net_),
            .in3(N__3051),
            .lcout(\row_counter.internal_count_9 ),
            .ltout(),
            .carryin(\row_counter.n751 ),
            .carryout(\row_counter.n752 ),
            .clk(N__3802),
            .ce(N__3437),
            .sr(N__3923));
    defparam \row_counter.internal_count__i10_LC_5_8_2 .C_ON=1'b1;
    defparam \row_counter.internal_count__i10_LC_5_8_2 .SEQ_MODE=4'b1000;
    defparam \row_counter.internal_count__i10_LC_5_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \row_counter.internal_count__i10_LC_5_8_2  (
            .in0(_gnd_net_),
            .in1(N__3723),
            .in2(_gnd_net_),
            .in3(N__3093),
            .lcout(\row_counter.internal_count_10 ),
            .ltout(),
            .carryin(\row_counter.n752 ),
            .carryout(\row_counter.n753 ),
            .clk(N__3802),
            .ce(N__3437),
            .sr(N__3923));
    defparam \row_counter.internal_count__i11_LC_5_8_3 .C_ON=1'b1;
    defparam \row_counter.internal_count__i11_LC_5_8_3 .SEQ_MODE=4'b1000;
    defparam \row_counter.internal_count__i11_LC_5_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \row_counter.internal_count__i11_LC_5_8_3  (
            .in0(_gnd_net_),
            .in1(N__3708),
            .in2(_gnd_net_),
            .in3(N__3090),
            .lcout(\row_counter.internal_count_11 ),
            .ltout(),
            .carryin(\row_counter.n753 ),
            .carryout(\row_counter.n754 ),
            .clk(N__3802),
            .ce(N__3437),
            .sr(N__3923));
    defparam \row_counter.internal_count__i12_LC_5_8_4 .C_ON=1'b1;
    defparam \row_counter.internal_count__i12_LC_5_8_4 .SEQ_MODE=4'b1000;
    defparam \row_counter.internal_count__i12_LC_5_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \row_counter.internal_count__i12_LC_5_8_4  (
            .in0(_gnd_net_),
            .in1(N__3693),
            .in2(_gnd_net_),
            .in3(N__3087),
            .lcout(\row_counter.internal_count_12 ),
            .ltout(),
            .carryin(\row_counter.n754 ),
            .carryout(\row_counter.n755 ),
            .clk(N__3802),
            .ce(N__3437),
            .sr(N__3923));
    defparam \row_counter.internal_count__i13_LC_5_8_5 .C_ON=1'b1;
    defparam \row_counter.internal_count__i13_LC_5_8_5 .SEQ_MODE=4'b1000;
    defparam \row_counter.internal_count__i13_LC_5_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \row_counter.internal_count__i13_LC_5_8_5  (
            .in0(_gnd_net_),
            .in1(N__3678),
            .in2(_gnd_net_),
            .in3(N__3084),
            .lcout(\row_counter.internal_count_13 ),
            .ltout(),
            .carryin(\row_counter.n755 ),
            .carryout(\row_counter.n756 ),
            .clk(N__3802),
            .ce(N__3437),
            .sr(N__3923));
    defparam \row_counter.internal_count__i14_LC_5_8_6 .C_ON=1'b1;
    defparam \row_counter.internal_count__i14_LC_5_8_6 .SEQ_MODE=4'b1000;
    defparam \row_counter.internal_count__i14_LC_5_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \row_counter.internal_count__i14_LC_5_8_6  (
            .in0(_gnd_net_),
            .in1(N__3663),
            .in2(_gnd_net_),
            .in3(N__3081),
            .lcout(\row_counter.internal_count_14 ),
            .ltout(),
            .carryin(\row_counter.n756 ),
            .carryout(\row_counter.n757 ),
            .clk(N__3802),
            .ce(N__3437),
            .sr(N__3923));
    defparam \row_counter.internal_count__i15_LC_5_8_7 .C_ON=1'b0;
    defparam \row_counter.internal_count__i15_LC_5_8_7 .SEQ_MODE=4'b1000;
    defparam \row_counter.internal_count__i15_LC_5_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \row_counter.internal_count__i15_LC_5_8_7  (
            .in0(_gnd_net_),
            .in1(N__3648),
            .in2(_gnd_net_),
            .in3(N__3078),
            .lcout(\row_counter.internal_count_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3802),
            .ce(N__3437),
            .sr(N__3923));
    defparam CONSTANT_ONE_LUT4_LC_5_9_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_5_9_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_5_9_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_5_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.output_enable_I_0_i1_2_lut_LC_5_9_4 .C_ON=1'b0;
    defparam \row_sr.output_enable_I_0_i1_2_lut_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \row_sr.output_enable_I_0_i1_2_lut_LC_5_9_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \row_sr.output_enable_I_0_i1_2_lut_LC_5_9_4  (
            .in0(N__3114),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4619),
            .lcout(sr_row_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.output_enable_I_0_i5_2_lut_LC_5_9_5 .C_ON=1'b0;
    defparam \row_sr.output_enable_I_0_i5_2_lut_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \row_sr.output_enable_I_0_i5_2_lut_LC_5_9_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \row_sr.output_enable_I_0_i5_2_lut_LC_5_9_5  (
            .in0(N__4620),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4416),
            .lcout(sr_row_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.output_enable_I_0_i8_2_lut_LC_5_9_6 .C_ON=1'b0;
    defparam \row_sr.output_enable_I_0_i8_2_lut_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \row_sr.output_enable_I_0_i8_2_lut_LC_5_9_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \row_sr.output_enable_I_0_i8_2_lut_LC_5_9_6  (
            .in0(_gnd_net_),
            .in1(N__4621),
            .in2(_gnd_net_),
            .in3(N__4320),
            .lcout(sr_row_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_7_LC_5_9_7.C_ON=1'b0;
    defparam i1_3_lut_adj_7_LC_5_9_7.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_7_LC_5_9_7.LUT_INIT=16'b1111111100100010;
    LogicCell40 i1_3_lut_adj_7_LC_5_9_7 (
            .in0(N__3456),
            .in1(N__3820),
            .in2(_gnd_net_),
            .in3(N__3913),
            .lcout(n189),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.shifted_data_i1_LC_5_10_2 .C_ON=1'b0;
    defparam \divider_sr.shifted_data_i1_LC_5_10_2 .SEQ_MODE=4'b1000;
    defparam \divider_sr.shifted_data_i1_LC_5_10_2 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \divider_sr.shifted_data_i1_LC_5_10_2  (
            .in0(N__3389),
            .in1(N__3318),
            .in2(N__3374),
            .in3(N__3242),
            .lcout(shifted_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4710),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.shifted_data_i0_LC_5_10_3 .C_ON=1'b0;
    defparam \divider_sr.shifted_data_i0_LC_5_10_3 .SEQ_MODE=4'b1000;
    defparam \divider_sr.shifted_data_i0_LC_5_10_3 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \divider_sr.shifted_data_i0_LC_5_10_3  (
            .in0(N__3317),
            .in1(N__3420),
            .in2(N__3248),
            .in3(N__3388),
            .lcout(shifted_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4710),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.shifted_data_i3_LC_5_10_4 .C_ON=1'b0;
    defparam \divider_sr.shifted_data_i3_LC_5_10_4 .SEQ_MODE=4'b1000;
    defparam \divider_sr.shifted_data_i3_LC_5_10_4 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \divider_sr.shifted_data_i3_LC_5_10_4  (
            .in0(N__3244),
            .in1(N__3343),
            .in2(N__3164),
            .in3(N__3320),
            .lcout(shifted_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4710),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.shifted_data_i2_LC_5_10_6 .C_ON=1'b0;
    defparam \divider_sr.shifted_data_i2_LC_5_10_6 .SEQ_MODE=4'b1000;
    defparam \divider_sr.shifted_data_i2_LC_5_10_6 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \divider_sr.shifted_data_i2_LC_5_10_6  (
            .in0(N__3243),
            .in1(N__3367),
            .in2(N__3351),
            .in3(N__3319),
            .lcout(shifted_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4710),
            .ce(),
            .sr(_gnd_net_));
    defparam \divider_sr.shifted_data_i4_LC_5_11_7 .C_ON=1'b0;
    defparam \divider_sr.shifted_data_i4_LC_5_11_7 .SEQ_MODE=4'b1000;
    defparam \divider_sr.shifted_data_i4_LC_5_11_7 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \divider_sr.shifted_data_i4_LC_5_11_7  (
            .in0(N__3324),
            .in1(N__3133),
            .in2(N__3252),
            .in3(N__3160),
            .lcout(shifted_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4712),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.shifted_data_i1_LC_6_6_2 .C_ON=1'b0;
    defparam \row_sr.shifted_data_i1_LC_6_6_2 .SEQ_MODE=4'b1000;
    defparam \row_sr.shifted_data_i1_LC_6_6_2 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \row_sr.shifted_data_i1_LC_6_6_2  (
            .in0(N__4965),
            .in1(N__3631),
            .in2(N__4879),
            .in3(N__3110),
            .lcout(shifted_data_1_adj_114),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4717),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.output_enable_I_0_i2_2_lut_LC_6_6_3 .C_ON=1'b0;
    defparam \row_sr.output_enable_I_0_i2_2_lut_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \row_sr.output_enable_I_0_i2_2_lut_LC_6_6_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \row_sr.output_enable_I_0_i2_2_lut_LC_6_6_3  (
            .in0(N__3633),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4645),
            .lcout(sr_row_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.shifted_data_i2_LC_6_6_4 .C_ON=1'b0;
    defparam \row_sr.shifted_data_i2_LC_6_6_4 .SEQ_MODE=4'b1000;
    defparam \row_sr.shifted_data_i2_LC_6_6_4 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \row_sr.shifted_data_i2_LC_6_6_4  (
            .in0(N__4966),
            .in1(N__4450),
            .in2(N__4880),
            .in3(N__3632),
            .lcout(shifted_data_2_adj_113),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4717),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_counter.sub_8_add_2_2_lut_LC_6_7_0 .C_ON=1'b1;
    defparam \row_counter.sub_8_add_2_2_lut_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \row_counter.sub_8_add_2_2_lut_LC_6_7_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \row_counter.sub_8_add_2_2_lut_LC_6_7_0  (
            .in0(N__3621),
            .in1(N__3609),
            .in2(_gnd_net_),
            .in3(N__3600),
            .lcout(n1),
            .ltout(),
            .carryin(bfn_6_7_0_),
            .carryout(\row_counter.n696 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_counter.sub_8_add_2_3_lut_LC_6_7_1 .C_ON=1'b1;
    defparam \row_counter.sub_8_add_2_3_lut_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \row_counter.sub_8_add_2_3_lut_LC_6_7_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \row_counter.sub_8_add_2_3_lut_LC_6_7_1  (
            .in0(N__3597),
            .in1(N__4120),
            .in2(N__3585),
            .in3(N__3576),
            .lcout(n2),
            .ltout(),
            .carryin(\row_counter.n696 ),
            .carryout(\row_counter.n697 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_counter.sub_8_add_2_4_lut_LC_6_7_2 .C_ON=1'b1;
    defparam \row_counter.sub_8_add_2_4_lut_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \row_counter.sub_8_add_2_4_lut_LC_6_7_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \row_counter.sub_8_add_2_4_lut_LC_6_7_2  (
            .in0(N__3572),
            .in1(N__4434),
            .in2(N__4143),
            .in3(N__3558),
            .lcout(n3),
            .ltout(),
            .carryin(\row_counter.n697 ),
            .carryout(\row_counter.n698 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_counter.sub_8_add_2_5_lut_LC_6_7_3 .C_ON=1'b1;
    defparam \row_counter.sub_8_add_2_5_lut_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \row_counter.sub_8_add_2_5_lut_LC_6_7_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \row_counter.sub_8_add_2_5_lut_LC_6_7_3  (
            .in0(N__3555),
            .in1(N__4124),
            .in2(N__4464),
            .in3(N__3540),
            .lcout(n4),
            .ltout(),
            .carryin(\row_counter.n698 ),
            .carryout(\row_counter.n699 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_counter.sub_8_add_2_6_lut_LC_6_7_4 .C_ON=1'b1;
    defparam \row_counter.sub_8_add_2_6_lut_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \row_counter.sub_8_add_2_6_lut_LC_6_7_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \row_counter.sub_8_add_2_6_lut_LC_6_7_4  (
            .in0(N__3536),
            .in1(N__3525),
            .in2(N__4144),
            .in3(N__3516),
            .lcout(n5),
            .ltout(),
            .carryin(\row_counter.n699 ),
            .carryout(\row_counter.n700 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_counter.sub_8_add_2_7_lut_LC_6_7_5 .C_ON=1'b1;
    defparam \row_counter.sub_8_add_2_7_lut_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \row_counter.sub_8_add_2_7_lut_LC_6_7_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \row_counter.sub_8_add_2_7_lut_LC_6_7_5  (
            .in0(N__3513),
            .in1(N__4128),
            .in2(N__4662),
            .in3(N__3501),
            .lcout(n6),
            .ltout(),
            .carryin(\row_counter.n700 ),
            .carryout(\row_counter.n701 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_counter.sub_8_add_2_8_lut_LC_6_7_6 .C_ON=1'b1;
    defparam \row_counter.sub_8_add_2_8_lut_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \row_counter.sub_8_add_2_8_lut_LC_6_7_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \row_counter.sub_8_add_2_8_lut_LC_6_7_6  (
            .in0(N__3497),
            .in1(N__4008),
            .in2(N__4145),
            .in3(N__3486),
            .lcout(n7_adj_121),
            .ltout(),
            .carryin(\row_counter.n701 ),
            .carryout(\row_counter.n702 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_counter.sub_8_add_2_9_lut_LC_6_7_7 .C_ON=1'b1;
    defparam \row_counter.sub_8_add_2_9_lut_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \row_counter.sub_8_add_2_9_lut_LC_6_7_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \row_counter.sub_8_add_2_9_lut_LC_6_7_7  (
            .in0(N__3482),
            .in1(N__4132),
            .in2(N__3471),
            .in3(N__3459),
            .lcout(n8_adj_122),
            .ltout(),
            .carryin(\row_counter.n702 ),
            .carryout(\row_counter.n703 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_counter.sub_8_add_2_10_lut_LC_6_8_0 .C_ON=1'b1;
    defparam \row_counter.sub_8_add_2_10_lut_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \row_counter.sub_8_add_2_10_lut_LC_6_8_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \row_counter.sub_8_add_2_10_lut_LC_6_8_0  (
            .in0(N__3755),
            .in1(N__4014),
            .in2(N__4111),
            .in3(N__3744),
            .lcout(n9_adj_123),
            .ltout(),
            .carryin(bfn_6_8_0_),
            .carryout(\row_counter.n704 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_counter.sub_8_add_2_11_lut_LC_6_8_1 .C_ON=1'b1;
    defparam \row_counter.sub_8_add_2_11_lut_LC_6_8_1 .SEQ_MODE=4'b0000;
    defparam \row_counter.sub_8_add_2_11_lut_LC_6_8_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \row_counter.sub_8_add_2_11_lut_LC_6_8_1  (
            .in0(N__3741),
            .in1(N__3999),
            .in2(N__4115),
            .in3(N__3726),
            .lcout(n10_adj_124),
            .ltout(),
            .carryin(\row_counter.n704 ),
            .carryout(\row_counter.n705 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_counter.sub_8_add_2_12_lut_LC_6_8_2 .C_ON=1'b1;
    defparam \row_counter.sub_8_add_2_12_lut_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \row_counter.sub_8_add_2_12_lut_LC_6_8_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \row_counter.sub_8_add_2_12_lut_LC_6_8_2  (
            .in0(N__3722),
            .in1(N__4236),
            .in2(N__4112),
            .in3(N__3711),
            .lcout(n11_adj_125),
            .ltout(),
            .carryin(\row_counter.n705 ),
            .carryout(\row_counter.n706 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_counter.sub_8_add_2_13_lut_LC_6_8_3 .C_ON=1'b1;
    defparam \row_counter.sub_8_add_2_13_lut_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \row_counter.sub_8_add_2_13_lut_LC_6_8_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \row_counter.sub_8_add_2_13_lut_LC_6_8_3  (
            .in0(N__3707),
            .in1(N__4287),
            .in2(N__4116),
            .in3(N__3696),
            .lcout(n12_adj_126),
            .ltout(),
            .carryin(\row_counter.n706 ),
            .carryout(\row_counter.n707 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_counter.sub_8_add_2_14_lut_LC_6_8_4 .C_ON=1'b1;
    defparam \row_counter.sub_8_add_2_14_lut_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \row_counter.sub_8_add_2_14_lut_LC_6_8_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \row_counter.sub_8_add_2_14_lut_LC_6_8_4  (
            .in0(N__3692),
            .in1(N__5034),
            .in2(N__4113),
            .in3(N__3681),
            .lcout(\row_counter.n13 ),
            .ltout(),
            .carryin(\row_counter.n707 ),
            .carryout(\row_counter.n708 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_counter.sub_8_add_2_15_lut_LC_6_8_5 .C_ON=1'b1;
    defparam \row_counter.sub_8_add_2_15_lut_LC_6_8_5 .SEQ_MODE=4'b0000;
    defparam \row_counter.sub_8_add_2_15_lut_LC_6_8_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \row_counter.sub_8_add_2_15_lut_LC_6_8_5  (
            .in0(N__3677),
            .in1(N__4269),
            .in2(N__4117),
            .in3(N__3666),
            .lcout(n14_adj_127),
            .ltout(),
            .carryin(\row_counter.n708 ),
            .carryout(\row_counter.n709 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_counter.sub_8_add_2_16_lut_LC_6_8_6 .C_ON=1'b1;
    defparam \row_counter.sub_8_add_2_16_lut_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \row_counter.sub_8_add_2_16_lut_LC_6_8_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \row_counter.sub_8_add_2_16_lut_LC_6_8_6  (
            .in0(N__3662),
            .in1(N__4296),
            .in2(N__4114),
            .in3(N__3651),
            .lcout(n15_adj_128),
            .ltout(),
            .carryin(\row_counter.n709 ),
            .carryout(\row_counter.n710 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_counter.sub_8_add_2_17_lut_LC_6_8_7 .C_ON=1'b1;
    defparam \row_counter.sub_8_add_2_17_lut_LC_6_8_7 .SEQ_MODE=4'b0000;
    defparam \row_counter.sub_8_add_2_17_lut_LC_6_8_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \row_counter.sub_8_add_2_17_lut_LC_6_8_7  (
            .in0(N__3647),
            .in1(N__4278),
            .in2(N__4118),
            .in3(N__3636),
            .lcout(n16_adj_129),
            .ltout(),
            .carryin(\row_counter.n710 ),
            .carryout(\row_counter.n711 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_counter.sub_8_add_2_18_lut_LC_6_9_0 .C_ON=1'b0;
    defparam \row_counter.sub_8_add_2_18_lut_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \row_counter.sub_8_add_2_18_lut_LC_6_9_0 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \row_counter.sub_8_add_2_18_lut_LC_6_9_0  (
            .in0(N__4227),
            .in1(N__4062),
            .in2(_gnd_net_),
            .in3(N__4017),
            .lcout(n775),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.output_enable_I_0_i9_2_lut_LC_6_9_1 .C_ON=1'b0;
    defparam \row_sr.output_enable_I_0_i9_2_lut_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \row_sr.output_enable_I_0_i9_2_lut_LC_6_9_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \row_sr.output_enable_I_0_i9_2_lut_LC_6_9_1  (
            .in0(N__4648),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5049),
            .lcout(sr_row_data_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.output_enable_I_0_i7_2_lut_LC_6_9_2 .C_ON=1'b0;
    defparam \row_sr.output_enable_I_0_i7_2_lut_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \row_sr.output_enable_I_0_i7_2_lut_LC_6_9_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \row_sr.output_enable_I_0_i7_2_lut_LC_6_9_2  (
            .in0(_gnd_net_),
            .in1(N__4647),
            .in2(_gnd_net_),
            .in3(N__4341),
            .lcout(sr_row_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.output_enable_I_0_i10_2_lut_LC_6_9_3 .C_ON=1'b0;
    defparam \row_sr.output_enable_I_0_i10_2_lut_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \row_sr.output_enable_I_0_i10_2_lut_LC_6_9_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \row_sr.output_enable_I_0_i10_2_lut_LC_6_9_3  (
            .in0(N__4646),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4754),
            .lcout(sr_row_data_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i748_2_lut_LC_6_9_4.C_ON=1'b0;
    defparam i748_2_lut_LC_6_9_4.SEQ_MODE=4'b0000;
    defparam i748_2_lut_LC_6_9_4.LUT_INIT=16'b1111111111001100;
    LogicCell40 i748_2_lut_LC_6_9_4 (
            .in0(_gnd_net_),
            .in1(N__3993),
            .in2(_gnd_net_),
            .in3(N__3984),
            .lcout(),
            .ltout(n811_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i768_4_lut_LC_6_9_5.C_ON=1'b0;
    defparam i768_4_lut_LC_6_9_5.SEQ_MODE=4'b0000;
    defparam i768_4_lut_LC_6_9_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i768_4_lut_LC_6_9_5 (
            .in0(N__3975),
            .in1(N__3966),
            .in2(N__3960),
            .in3(N__3957),
            .lcout(),
            .ltout(n831_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i772_4_lut_LC_6_9_6.C_ON=1'b0;
    defparam i772_4_lut_LC_6_9_6.SEQ_MODE=4'b0000;
    defparam i772_4_lut_LC_6_9_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i772_4_lut_LC_6_9_6 (
            .in0(N__3948),
            .in1(N__3939),
            .in2(N__3933),
            .in3(N__3930),
            .lcout(),
            .ltout(n835_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_counter.internal_count_reached_18_LC_6_9_7 .C_ON=1'b0;
    defparam \row_counter.internal_count_reached_18_LC_6_9_7 .SEQ_MODE=4'b1000;
    defparam \row_counter.internal_count_reached_18_LC_6_9_7 .LUT_INIT=16'b0010001000100011;
    LogicCell40 \row_counter.internal_count_reached_18_LC_6_9_7  (
            .in0(N__3821),
            .in1(N__3914),
            .in2(N__3831),
            .in3(N__4347),
            .lcout(row_complete),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3804),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.output_enable_I_0_i15_2_lut_LC_6_10_0 .C_ON=1'b0;
    defparam \row_sr.output_enable_I_0_i15_2_lut_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \row_sr.output_enable_I_0_i15_2_lut_LC_6_10_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \row_sr.output_enable_I_0_i15_2_lut_LC_6_10_0  (
            .in0(N__4630),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4248),
            .lcout(sr_row_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.output_enable_I_0_i12_2_lut_LC_6_10_1 .C_ON=1'b0;
    defparam \row_sr.output_enable_I_0_i12_2_lut_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \row_sr.output_enable_I_0_i12_2_lut_LC_6_10_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \row_sr.output_enable_I_0_i12_2_lut_LC_6_10_1  (
            .in0(N__5003),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4628),
            .lcout(sr_row_data_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.shifted_data_i11_LC_6_10_2 .C_ON=1'b0;
    defparam \row_sr.shifted_data_i11_LC_6_10_2 .SEQ_MODE=4'b1000;
    defparam \row_sr.shifted_data_i11_LC_6_10_2 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \row_sr.shifted_data_i11_LC_6_10_2  (
            .in0(N__4961),
            .in1(N__5002),
            .in2(N__4862),
            .in3(N__4733),
            .lcout(shifted_data_11_adj_104),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4711),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.output_enable_I_0_i16_2_lut_LC_6_10_3 .C_ON=1'b0;
    defparam \row_sr.output_enable_I_0_i16_2_lut_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \row_sr.output_enable_I_0_i16_2_lut_LC_6_10_3 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \row_sr.output_enable_I_0_i16_2_lut_LC_6_10_3  (
            .in0(N__4259),
            .in1(N__4631),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sr_row_data_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.output_enable_I_0_i14_2_lut_LC_6_10_4 .C_ON=1'b0;
    defparam \row_sr.output_enable_I_0_i14_2_lut_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \row_sr.output_enable_I_0_i14_2_lut_LC_6_10_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \row_sr.output_enable_I_0_i14_2_lut_LC_6_10_4  (
            .in0(N__4629),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5024),
            .lcout(sr_row_data_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.shifted_data_i15_LC_6_10_5 .C_ON=1'b0;
    defparam \row_sr.shifted_data_i15_LC_6_10_5 .SEQ_MODE=4'b1000;
    defparam \row_sr.shifted_data_i15_LC_6_10_5 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \row_sr.shifted_data_i15_LC_6_10_5  (
            .in0(N__4247),
            .in1(N__4963),
            .in2(N__4260),
            .in3(N__4835),
            .lcout(shifted_data_15_adj_100),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4711),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.shifted_data_i14_LC_6_10_6 .C_ON=1'b0;
    defparam \row_sr.shifted_data_i14_LC_6_10_6 .SEQ_MODE=4'b1000;
    defparam \row_sr.shifted_data_i14_LC_6_10_6 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \row_sr.shifted_data_i14_LC_6_10_6  (
            .in0(N__4962),
            .in1(N__4246),
            .in2(N__4863),
            .in3(N__5023),
            .lcout(shifted_data_14_adj_101),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4711),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.output_enable_I_0_i11_2_lut_LC_6_10_7 .C_ON=1'b0;
    defparam \row_sr.output_enable_I_0_i11_2_lut_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \row_sr.output_enable_I_0_i11_2_lut_LC_6_10_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \row_sr.output_enable_I_0_i11_2_lut_LC_6_10_7  (
            .in0(N__4734),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4627),
            .lcout(sr_row_data_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.shifted_data_i3_LC_7_6_0 .C_ON=1'b0;
    defparam \row_sr.shifted_data_i3_LC_7_6_0 .SEQ_MODE=4'b1000;
    defparam \row_sr.shifted_data_i3_LC_7_6_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \row_sr.shifted_data_i3_LC_7_6_0  (
            .in0(N__4976),
            .in1(N__4480),
            .in2(N__4877),
            .in3(N__4451),
            .lcout(shifted_data_3_adj_112),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4719),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.shifted_data_i5_LC_7_7_0 .C_ON=1'b0;
    defparam \row_sr.shifted_data_i5_LC_7_7_0 .SEQ_MODE=4'b1000;
    defparam \row_sr.shifted_data_i5_LC_7_7_0 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \row_sr.shifted_data_i5_LC_7_7_0  (
            .in0(N__4408),
            .in1(N__4872),
            .in2(N__4977),
            .in3(N__4675),
            .lcout(shifted_data_5_adj_110),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4718),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.output_enable_I_0_i3_2_lut_LC_7_7_2 .C_ON=1'b0;
    defparam \row_sr.output_enable_I_0_i3_2_lut_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \row_sr.output_enable_I_0_i3_2_lut_LC_7_7_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \row_sr.output_enable_I_0_i3_2_lut_LC_7_7_2  (
            .in0(N__4650),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4452),
            .lcout(sr_row_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i740_2_lut_LC_7_7_4.C_ON=1'b0;
    defparam i740_2_lut_LC_7_7_4.SEQ_MODE=4'b0000;
    defparam i740_2_lut_LC_7_7_4.LUT_INIT=16'b1111111111001100;
    LogicCell40 i740_2_lut_LC_7_7_4 (
            .in0(_gnd_net_),
            .in1(N__4428),
            .in2(_gnd_net_),
            .in3(N__4422),
            .lcout(n803),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.shifted_data_i6_LC_7_7_5 .C_ON=1'b0;
    defparam \row_sr.shifted_data_i6_LC_7_7_5 .SEQ_MODE=4'b1000;
    defparam \row_sr.shifted_data_i6_LC_7_7_5 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \row_sr.shifted_data_i6_LC_7_7_5  (
            .in0(N__4676),
            .in1(N__4975),
            .in2(N__4881),
            .in3(N__4336),
            .lcout(shifted_data_6_adj_109),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4718),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.shifted_data_i4_LC_7_7_7 .C_ON=1'b0;
    defparam \row_sr.shifted_data_i4_LC_7_7_7 .SEQ_MODE=4'b1000;
    defparam \row_sr.shifted_data_i4_LC_7_7_7 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \row_sr.shifted_data_i4_LC_7_7_7  (
            .in0(N__4871),
            .in1(N__4971),
            .in2(N__4488),
            .in3(N__4409),
            .lcout(shifted_data_4_adj_111),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4718),
            .ce(),
            .sr(_gnd_net_));
    defparam i730_4_lut_LC_7_8_2.C_ON=1'b0;
    defparam i730_4_lut_LC_7_8_2.SEQ_MODE=4'b0000;
    defparam i730_4_lut_LC_7_8_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i730_4_lut_LC_7_8_2 (
            .in0(N__4395),
            .in1(N__4389),
            .in2(N__4383),
            .in3(N__4374),
            .lcout(),
            .ltout(n793_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i766_4_lut_LC_7_8_3.C_ON=1'b0;
    defparam i766_4_lut_LC_7_8_3.SEQ_MODE=4'b0000;
    defparam i766_4_lut_LC_7_8_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i766_4_lut_LC_7_8_3 (
            .in0(N__4368),
            .in1(N__4362),
            .in2(N__4356),
            .in3(N__4353),
            .lcout(n829),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.shifted_data_i7_LC_7_8_5 .C_ON=1'b0;
    defparam \row_sr.shifted_data_i7_LC_7_8_5 .SEQ_MODE=4'b1000;
    defparam \row_sr.shifted_data_i7_LC_7_8_5 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \row_sr.shifted_data_i7_LC_7_8_5  (
            .in0(N__4970),
            .in1(N__4312),
            .in2(N__4876),
            .in3(N__4337),
            .lcout(shifted_data_7_adj_108),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4715),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.shifted_data_i8_LC_7_9_0 .C_ON=1'b0;
    defparam \row_sr.shifted_data_i8_LC_7_9_0 .SEQ_MODE=4'b1000;
    defparam \row_sr.shifted_data_i8_LC_7_9_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \row_sr.shifted_data_i8_LC_7_9_0  (
            .in0(N__4924),
            .in1(N__5047),
            .in2(N__4828),
            .in3(N__4313),
            .lcout(shifted_data_8_adj_107),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4714),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.shifted_data_i9_LC_7_9_7 .C_ON=1'b0;
    defparam \row_sr.shifted_data_i9_LC_7_9_7 .SEQ_MODE=4'b1000;
    defparam \row_sr.shifted_data_i9_LC_7_9_7 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \row_sr.shifted_data_i9_LC_7_9_7  (
            .in0(N__5048),
            .in1(N__4798),
            .in2(N__4755),
            .in3(N__4925),
            .lcout(shifted_data_9_adj_106),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4714),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.output_enable_I_0_i13_2_lut_LC_7_10_1 .C_ON=1'b0;
    defparam \row_sr.output_enable_I_0_i13_2_lut_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \row_sr.output_enable_I_0_i13_2_lut_LC_7_10_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \row_sr.output_enable_I_0_i13_2_lut_LC_7_10_1  (
            .in0(N__4649),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4989),
            .lcout(sr_row_data_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.shifted_data_i13_LC_7_10_3 .C_ON=1'b0;
    defparam \row_sr.shifted_data_i13_LC_7_10_3 .SEQ_MODE=4'b1000;
    defparam \row_sr.shifted_data_i13_LC_7_10_3 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \row_sr.shifted_data_i13_LC_7_10_3  (
            .in0(N__4840),
            .in1(N__4988),
            .in2(N__5025),
            .in3(N__4969),
            .lcout(shifted_data_13_adj_102),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4713),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.shifted_data_i12_LC_7_10_5 .C_ON=1'b0;
    defparam \row_sr.shifted_data_i12_LC_7_10_5 .SEQ_MODE=4'b1000;
    defparam \row_sr.shifted_data_i12_LC_7_10_5 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \row_sr.shifted_data_i12_LC_7_10_5  (
            .in0(N__4839),
            .in1(N__4987),
            .in2(N__5007),
            .in3(N__4968),
            .lcout(shifted_data_12_adj_103),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4713),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.shifted_data_i10_LC_7_10_6 .C_ON=1'b0;
    defparam \row_sr.shifted_data_i10_LC_7_10_6 .SEQ_MODE=4'b1000;
    defparam \row_sr.shifted_data_i10_LC_7_10_6 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \row_sr.shifted_data_i10_LC_7_10_6  (
            .in0(N__4967),
            .in1(N__4732),
            .in2(N__4864),
            .in3(N__4753),
            .lcout(shifted_data_10_adj_105),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4713),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.output_enable_I_0_i6_2_lut_LC_8_7_1 .C_ON=1'b0;
    defparam \row_sr.output_enable_I_0_i6_2_lut_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \row_sr.output_enable_I_0_i6_2_lut_LC_8_7_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \row_sr.output_enable_I_0_i6_2_lut_LC_8_7_1  (
            .in0(N__4677),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4544),
            .lcout(sr_row_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \row_sr.output_enable_I_0_i4_2_lut_LC_8_7_4 .C_ON=1'b0;
    defparam \row_sr.output_enable_I_0_i4_2_lut_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \row_sr.output_enable_I_0_i4_2_lut_LC_8_7_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \row_sr.output_enable_I_0_i4_2_lut_LC_8_7_4  (
            .in0(N__4543),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4484),
            .lcout(sr_row_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // top
